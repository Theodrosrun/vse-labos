`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
GNCxYQATjbMhzIJpeYg65fPHjq6uKtdDkmMi2LWymXyvg+oN2+wQzONkmYD6HUv8
QTeesv95Cxz3s+G58OqDGvK6UvRoIbUTeTXNZ7wnF6aJjtOkf72DAcT3KWTb+PCL
blDoPBv+GvOkz5QEzMQXguXzDhitpe4/3jWP/X0Ic6YYV90lJ77O2Gvk7kC1x4Fw
8nJVQaiiihcANnY+fgyLnJQ4hP/lfes8Kg9TfrHtG1okzIqxBfeQOK5emnMyVoLc
eg2eUki+4gQ6fbmoH6vSYqTCdjVmWJbd+7ZNrLofbfqt8fcPM3F/ds3/qZC/oNp6
m5uhaAMKpMbOAP1xRWjqbg==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5072 )
`protect data_block
RQ6vwd2Qewpp/E+FC2okyxtKdZzE+RhrM5oHxP0X9hbqVkeg3amRq7/y3TtDVk5F
DTvVggnAnvV3P13KOvohw3BObGTxcPCId9X8WeWryRzlHP6KxNSo2O4C/Takak7p
S82zyiuL/AzYz8d0/VDC1YscZt80EVgUIcUoTychsmbcWPgm34uTTmJ+dgUIskGT
+KzGcf/cT8R4yCrA99ZSs00xrcUXDLEwYRsexrHuMFEHBR4vrylM5FzFOXc7XYTl
Ql6HfXz2qLkIXdspDFFDR1nDBGlesw1XLGyFIfBBYFJFHTgPC3UAcdZlIcuYXsan
ZrknLsRvp3UhUq1MsBqU7xBsWPbDE9XAM2Vqh/tHTafBLp68ms9/ehSY8IMZjs+v
VbROfWnI5KV8XFXBk3AvH95mfIlNb8bNv/oA74yYNDGy6ZA3KJaWQNgAt/K0MaIP
kPjyVbZC4WKPSbEG8wzSdeJySkBGyfBFRYuxnBJnaMfKflgQlW7KR5+ArjDxi3p+
YtM4tIKblLh3sG52L1HOw1F+EQg6yJBkW5LWook/P4iZSGhlC3dagFCH2WkaASPi
he5GuvCFtaQExwzjnsLYtqMXGjU2tUWZSHpahNuvSB1P/bgwowck+ZjzG3yswvSO
r2HNi3iyMD47bx4SZSyAIYMgbeCU6UkLj8WJPCR9ciWE2Yx5CtGIUUruYtzrPmoY
aLiXKuC5tlXEqOzVZdKBe+YIxYtQlb2YTxuL4HrllFytVkBTa8oocSbOWhwWO90u
pSs94S1B3zFvkTSjra3dUVaWklpA+K8gwXu2nlS2yfpmpjRlAc4IpLsGla2XjzOT
A0fczL4VgrwCGNXj3VWUMrvUlRzICPbn/lNmFjpxWjSlIkHshnptDzqMIOmGnLs9
/w31Z+pfS5NRjgrXKZoV9O1c3OmMTDABsnrE/uO1s1NYItS5gub7bOfgPUEafmey
BILhyzuT8vnYllZ5Ivmaw97wkJkIF/IQQY3wBl54sZWpwc38R7TBc3KYVcNgpCGT
lRiTaoAgodFJkL8sCC2WPfeJAEe2GaOdvnmzcb+INxzSBjiPfSa5qMz2pKwVCTMe
SKs1Zs8nMPau9/xeEI6B28q3+3DSYZs5DHlVQ3XF0J2dfgSAm2yCzTULHg9VLQjV
xPwJzyiuHJ9hQCg5Iyve9mzECqyxQG7z7u5Ec08WHjVP0/Du6HYsE0yxsnj5lUQ2
RQ0HjBZkRdbkqAaBsIV2SQ59fTW2B+6ZzsHDIaKf5OTC97KHvp1ke4j8RJG4NY09
8HksS3vT2jeHRwUFDdJzXpqXcfDsdgN2cc6I3LC3vcgfA5Dzg4MewPgHvQtkRJhy
Qqt/gJQqEi0FgsRdqGho+soI6YzDcfUVD3+1ZTDz3GCKOx1dqvURdzgkdQ9o5Ks1
ykd/eEb2/gBCmwAGL15OrId+H02CkOgDe0E+hy3RKYMOZXX4pBlVZUehLzKiLxvW
gA5MNanq7TVuc51G2jFYCmn1hdKW4nMnRMjy+z6sY0A8xsfEpJksC32hH3bWLBGq
f2mN5DGPZZkX73nPxqDhmtuLapM3sl8WY2qbN1Nra3EvDwWwF6bWgwVaM0UY4tAi
JgX/jdLk5aMVxsmhnaVubLq3mvKcTf7zmiuL52HJnDL42O5v8zPtzcQtH/XXIQn5
QwdWWq0kqiasZ/tex6rD7ILb7bKMDKPUD6UhnNK9AgFmeF4zqFpUEXzVSQhARW7i
pmkQgm7nWS0UqWR6PicMcmUfHi9iImeXIZomoU4A7CkcBSMpKeD+18WsJ3rOFvZl
JZ36thxtEAijKp7CH14poMcA0QeEye7+ycCdG7rh7JWnjZf6lqwtd6kfKAB4BQYF
JArXHmyeMAc/UW+VoWwo6EC+fbPpqcNxOihx6mdLnagPz+7cnsTlUmTivylPEQWM
T7gd1Udl1M0eup1SI9Q5zRllymYQ8Mz++82t9lzJQXlg4M8Wr52/+wHBOLqVC/+t
B+fTjGufovj0uDvuDHjjl9fqigDAphuZ+Qvq/ghtkymp9+eVs2X/p3V6fNtS1Mxz
7hh3nhQHJ9xZDJhFssj1mcmuq5R+MxhPOiY2EPEiilgt4tGhfdc/tZ7QlMWBx02d
FTbNO4IfvD2ecAnHW1mRfsCoC13LZB0Nrt3GkW1YdCMUYrpPYju/dU5nvNYSuSIB
SStFw/C8bENyTMn9HDuXcJTktU9LANMpvumFDQlm7HLOmuhjkfB+B/d3gwm8/HI0
Jgw3U8+km0aBwkr5QVL1eUYucJL8CaVYMPepGTVtWQ329RLVmUQjNA9JnfE3J/TC
eDSrarrMLjfTGK9mNNaOL9ZG5IDulmRo/mV/l74L7hCw9hiKLfBXTFG2ezMkSazH
JvcmbTvW7Uj00DPRrGSVO/nepggAIRwfYnAEZ7Mgt+0PZf5arIxpgiPwb5n9tMjt
Ivp1037uGrU1pl2mpmwXQ4fqJ5kbWrSqvM8dsbwei3CjmdTxnhDysWDmlmiFKNpJ
xQqdX3qd4aJh6JDy4jIJWho3wPi/lYhfVdwk+EKmPGwVeoQSrPTbdZuzKPQjzEOz
hsSWn2RYD1WhSatRxje6DK4KnGB9d4hT7+cjFsSJK/YSsl2TC+HOkXgkLQfIGqSv
j4qIyC327ZqCBHw/uxke206fGuA3UKxs/KgPG7jCfwRenQwmWZ3PCGMcKr2+AgDT
ukspRaXrFPCEl3xp37zEiheZ/WceGj4My5m1ccLU0j38Rd8zzA4kPArt3Jms7m+q
s6insqppJ7pARg6CFuG48+0v+u31DeaClFS0qRYeMfW/oo1SQ/KCfCoHtAi0FjWf
A+1GwFZ8PnVFsOixfI0LFgn1G6qwzaSYBF1L14cr6NKSHz7+12lFruzBKN++gjq4
joGWLsAhzUbVtnkcqqUXZ7hrw52i8uY8HMo3Kv04XJCDR5SUsJjYpI8/H71vXue0
nuQjgFeMUjfseyJj0kAp9aH79NbGmV+Hzkt8G/9MjJbKMxkT3A/eOi/X4myA+aPK
S7nqclUVZG4wFDu3MtclkgzyW9ekri7c5Bs9oHjW/ZjgHCZYqLGUq1lUqXVejG/v
uNEshuIQwqoGAd7Hb0aIOjAPQeIOvyQMvUC6cKj68JCoQ2cRtPdgzlI4H9AY+sSL
pS1R8WSH2tz14ddJtr6gf83eS94ZsYUiw8++d1VdFvIDQjWMN2A+hXeZAnsLQfdZ
fObuJiLeqSroGI2yXFKskaBs6puk3e5GL40X05KYfC0fPj9cUie6RAeIlDaQ4dX6
QsH9jHj91xG5aFZyiv9ImATSlYw9mLeXg/FmdiK+t2VHMhwQ48Hp/pcDvDaCv8nw
7nI3RMHk7fVp+H+B0ATE/nylxxTZSmqhkC89v8WC8pLCr5e4p5xgYan2eHITDTnf
KaY5mgCEtjzO7wINAPc2abXgFlgpJ82RcXROqAwaHtJzcJ2572gfl6Zx7CUFJxBE
mgAd9HmVWiJQRtN2kPDCi05vKdFEcraTxZ2NLf4yAp781iwr7mvfRL65J5TY/a0v
xBLZj9TJlX1PtCJ0e9HEkVrTrVgPzSu06URZ0MqN6hw/jlAFiirUapd2Xu70NNz1
YHSE4kVpx514VgRriSN9OMbS8KRh6JECVHp4kMwvk0uTFPpN+OQNOMGCgXIAJnXA
RIJLRIszmNMBlIfrAp0ALc3tF1In87A7eKPzQgkQ8ytVUBLcwxrzbH9JN8ml7AyW
Lh9Bnn2VaYOcmeKfjkLMi8hXI0DZvZ1uxd6Np/5dAnr5ptCXX0BHUKx0lVVACUWA
Ks/CSs8kCywecrcwRGjdb5UCAis/bkXOdotheB1XHCd3ZW0NpBe+Zzr47+mC845f
+QTCYaaKzJ+dN6AB1amsGwSLt47zZL5PV66x0+TdN/ghueSvyvvq6B1iqgK0sW0J
x8Estt6VBfbsJ1REHiOh0vsBuMT6rA6Uc1o9xuBh6eOkbQMuyJv5vZf8aJux6H06
2a9XXEbBSsfBsLR1uwUbKrKYlje9tI536jOoyQ50R7aBb8lv8HGQOdDYjiYGPegy
7SKUUAqwKQRZWHlMUM2PCS+J2dhRQUHInQymuUnt8rmE6I7N5Bh6AapyZM5mxhGa
dPQI6MMkCyJV/Qjz4gbrC01vkhzL97yz3GStvCIysc26GpzYXVAAMvfytMdEAGjp
pM09XGqIvtq82oacTZkoOzXJ0Gp4HKl3bePaVHwGSk0kFG5SbsAGPeZHxRQeWOa2
chJUxDOgjoNupAFq7wMHEtQkpfdUTsUgPO+BOX01/OfoZoh5sSXEt6jkUAzTiV7e
DYBictR3uGaV1mZd3hduHr6e8Jbal+AB015fQZdIlfbCwQbsWyCmjhkYsuNmH3Wy
UD6pUkF3AQxmrLMh6QeMrAmFVZrjX7jgDhfsaEbBJtbPDO5RR3nOzgThHNX5nIpz
hqq+CCQjCxkK4u70awIxyRLOEy+NyMueH2YiCScKvkfGyA6eQ6gmRbML5YuPOyfT
Qz4Rwup7miigdwZfl+Y/JB/kXTS5QnSYBGDfHHEfbtzpXBB3o9Ug6DH7ZW2B89dB
B6ssezDUuLgiIR6KJKevFKNUjC5D4GdwlV5mo9OV1qDYPALM0w8+0CrApDxxsZEd
dxc9NXNXDTehaZxKr2Xdd/bEfvkllTAeUlTRoN1LhZ196s7XH+s0u4gL50fOS6ML
VMEwrRdIXznqknVYASuOcoSO5GM+hJV5RVM2d41fDMjnwpKS1w4PcVgQe4RSOcty
KmgYz5tCWm1WBRmeuAmlIjukv8g44CMMaqffD2CXf3acmd+tHCYJfbm/z3u8NtJw
4EHz4BS+TZ20xgkIjxKOAaBHn5qAr0fJwlhtGjLgM8VIEKoRrISF5B2iKvpKHDG2
xq2ZZsVury9PaG5X/YIYcSgp6d5Wf9GpropNdDKyYRmPzP+UkRcjaamzYWFwX7WP
UZrVeTih1IgFK/DxPDfff+BK1hu2xFfIKgmSh0MGR7n8U6yCSR2GHC4zVZDE27eM
6fkMiKBj9xE9ObDXGtWbJTOCuTuyTjfBhwu3B+DH4cbKKhLckkkGI5G2DSW+TpWJ
R8GhyWw9RfqFQniMp3tEQEUPbGAUzlrtRcZEwzWPQh/vHoxWv/UPdQDcfnR9ZkD1
uXs1H4jUOaI1aCRIhvzN8DU2b/HfjPCShdoDXWX5IvVCh7FDBsHgc7g38lM7hfqX
pZYD/JhcOnKBMhZ4w0J6n7FTzHBf35bPZbRBWuTbhOko4lRrymGe9g60/vxz0H/P
s8JbTbOlkytdFLrDuowkIFR/h8ncL3buzlQmNjgn39viaQDlF5K8qMlIBwOhLkd1
yqnA/jRrSf+jB/0LHYT76wMjX3MM7M783DTd03ZfdQJjgnksq67/5Ji+1GcVWRKb
6H0OaRnhF+rogxvm/ieIhQIVXTGrhrZ31TQp/yueW5XhcwN9/mkGBZE8BMslA2t9
UFxBBOmmufio9i8lvbPANANnufqb1J5ZughUDfTup7dGFjMBDu/Ruyr9mFi1P709
/uoFP8sYErshHO/2xc50hUl9jASY4xE74jIGG445EoZAL2f7+W0StgQZN7RhQbmB
wiv0sMtVlLT9lh0PYdxOYFDbjr81wV8vpz9+h6P5AbStiyb5T9a0SzFPJfO8QMGh
cHJ8Lv0UaDXE7Xct0Bl0DakXAEYU2P3tLMF8nLsYbqNFrcQL4JwQVyzgVW6qf+yj
ysRwwbqGniSnr2CtykcgYRV8Xqszf3mFpSdqOomu/p9DFtfZVKbeswnkJEllBnec
zuVbFP9vztvOVm/fjr6MMwFfN8rP9eH7rGwd/bAEqhdDoHmtE0WUD6xqSV6gL3Mn
6gKOKGbL47y4d+ruuCS7aHYGxzsriJH0kO9sb4Ea1tpDu9g2Sx737cMZb4BpgrX8
SFp3WAVUbR/yRjLQ+lpOpKwfKxVYb5t8rZt5qRj2CuhDlm14TLnKBO7hYPnrdO4S
4kWZ3I/cYlckh/wAYyvpkX5AQvDKEQJRGcWLOgEYUxUQ2bXt3DJpT12K522q55JJ
MBbjgOba/srMrw8AnOVXPi5JdHOy/FqW3Old8RJgpW6uWoQY7lRGw1Kgnhee4A9A
5XaCM6Q2Bevvg3LTkNEPufy9te3asmDc7JNUQ2jBWFwMLdHjcKjn8VKy+A/MvmB2
hJ7/cKE3uVS3rWMDP9qym2IZk+DarnJRdsPUl2MQTJ7DNnrCgnxuussn2FustWIB
hK1LxlOYugGICVoq7saWsJ1pbOUYMXHyB/WUluri/SfShjZo/oLnpBEuLvWZeOJW
MtRQf3AMV6PZP1/QjAelMPU6Hh4EJNmmc2vnrwcBAXblAvmsmA92Y4EnwA0sn4iR
vGAF5lgWmVH2H2j1Od6veInDdT3/VcbKdes7Q59jbiuDaQK8hwBwAn8gTJQ/MLqt
HzMKJ35UUnrKXg4XNbGHK9XACm1XlGrHVanfoC8uouMCfMnbworm0x2FiCFHfNDJ
wuBzE3Y0qeol4MXxRfd4MICu6iDgCyRd9sYg+oYz13w5iilNl0nlkUUt+dyfs3bX
7LDTEnuRU7+i+xk2oWtkqCDItUSTAQQ6pwrY0ZAREI1HBJBL87p461BUfM93/wsy
tyVpr/pGbR1wLQOtSWazHYyCv6NU0xv9Z9wQni+ib7YMUr8mu3y8MuOS0AfEBpMv
62MNx09saI4GitkZkBYOjwS/U4MQAIMSILaolpIy/QkBsDgoPbMfipZKKkwwrbud
ZKulMZIfKKuGqiy4pj0oaiyzkLlk5AaJX9xpQgbYh5A=
`protect end_protected
