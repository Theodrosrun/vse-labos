`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
jaadDojbPIt7kaASMldtDkOwWwZ4irMHQYp2GxAueXiUXhIsSAKrkWO4VEx+Byam
V4uIs5X56zM210+6dkPDe0Jg7gvJXM/mw7yPjsubaVZONhyOi2EmHbrskeZgS/qo
dGy7Y9eB1jkF4OMRcAUbybmCW8CWQNqkfSOZQcik1PV/P/xXktwqHZ5MYmhU7Fy+
FcS3vfDg/WE0zkjhXvnwMEFP2namwD/LFJdE55gUYKydK/eqdnSlEOMW0vmZAEjt
6V0Y8pD6qxcLxR2FUJK9+ary20xg3Wv5R5Wxy/4PS1xS+9oCeUdwtQ5h82Z92dgp
TRX2BygUptWtCdBO2vbpLA==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 28592 )
`protect data_block
ludPPAvlVCAFPgc1mGXaVMFrAOiT1ISeLUAs3j6mMSt302jZDbVPJK7nf+w2oerg
YWqklCikjPxKx+A8UYUWMacUcgKshQPxo5nzKibT8pknyUomjm4YcNHzEJK1pVbQ
ATTzJrIilZffyRdS8HkdzEzoiDWqvjPMS/pH+aiPCsk8f7JgvNJqxk2v7lCesWJ/
EHPs7yg/ssnBl7DsmXtKy3Km/B3SJ13e8dQ2mQ1ti25j6PK6Q1zQ34DmJZeB9TfA
6xzyQf2qQbWIpO4rW4klcAW0k2h6+irpMd1oh3DK1NGCKFUXNDo50cb6RzwS+x8D
lHE5BEDnMRbHft7eVQrow/CrPT+d8iaSO7NQccKM4K0QBJwc/dkIvMniBuhzpSOa
rTlophFssH7V9gJe7L6Uf3sM3Mg4uYZr2KuMABLM+nQmy4fIZqWl3Ec7tfwMody7
L6T3auGarlFajq2mUGYwN9975DmwAnxz2hlJmKkGegXpMOHf5k8iKxFYcx3muxoY
dkwpYVTNaYf2MCPYCA6BFgZmJCMOzSo57P0wpeNuCAap+6gjFaQT3i2StT7vNLRp
TJZxA4ZIC3hAwhJF6jGN6LU7dVgWsB8ZBSfqq7g8CQV4el/sWzaTRDqTsyhUeTLg
d0AIJ7M0j6bdURKPgTonhd3GTGzMXnoCZooSmIpaN9rR1TgF6sqPhPdPP958yHlZ
hxlKEPjCGLntdEnOaVkylj2vlVs+E2XSccVPxTu6vEApL9B6khfy6oOOt+5bUD7J
ruHOyvsQtPAVxSc7VAWsOB1LBNM08DPe3aYfI84kPVkAlZ+RPjO0b6WGq8JpgboG
BHptsNFc6/QYS0zjL6FJuJCUjNoJAzd/+y/UjWWCefsXPLaixOReFXiPK+7Jb3Jd
fMnvvjZSFdmFKBlFSfO4pGRvJgCwfnx9mGR20jojdi2w9xzbn1qtTt4D+KyjsIP4
3VeryYQrXKsvlPotyyv2fOXTto/IomBqLCD6Q2biehuZe3ppfxsItE60po0n6Zc2
2GmgrdgFG9TDxjB2imlKzzC0CSAaBEQAl5w46AL2AFlIFYb8u5Ngfk0cp+8+ZIUX
Wa5P1b4BKbYDCxZ26skaV16w/65tHcCwqN5LRppqL0fOjJKYEymInebSKDK/czuJ
L8oJ0bJ/YMlHR6UFMPpuoUEYOWgnP+pqTfsnyBC/W/PbcTo0u6C14Vee568FkE1V
tL1+fFPUnZKeDy6WD+96SHpF3xMbK7UmOc2KCi+1tOSjeHJKYvlSwJNWzPxW9hSo
ewXtM9HtAgPNOF6I3z3JvjMsZixLZBf1gZrMUQtcwTcM7Ul65+AZuSKId427Q8vO
5h6oS9cBxaKy5SywM0jaY0+n+YD3thhDjbr/j7e2wsx9ZFlGoXqcD76Foo/BUSrB
Pfjca0IsO8jJOsLmFDdm6lnk6vIYf7G0EnYoffdEb0l+ECdfiQVq6y2F/ih3G5zL
NswICxSK4/RMywDPgok3+vDFSCLfs59b4XH0x0fDozMdAwY0THL6ExGH0S0FYezI
QYdRAJJoVy/iFl0U2VYtMqGAZlOE4Fdvnyzn6ei6Ns19dz4Rcoa6Yfw60sOQuPPL
tmnU7QEw3MoQPiNxM1dHRg6U8n33s+U0wp7DStTdrndaDFZt20pSkRYKtKUjOY3Z
Zi2ZpPDecxHW3OVSO8uybqiCKaYwZDpfuoH2QqTqgfKxBnHwBJkCWBSXKPRSmVO1
fksi6gIQUfLrNHCgTnuacZzl/4dWmZLb6Z0/GWGfF5xlmSU7SGVFjIl0WZVBi6Kd
q5RapclnbD0tsKh3WU7uYxobZCh/IpOczqPsdkntESjk9yWc8J4FsPOdexN31NXJ
VL+YNBWVfN1hv+YCuLKvSEHvFCPme64oM7p8IqAj8DqXG2HTLgC+dKk1v3VERz5F
orbOstWCupdqr+rQ+RmxSj+gn74mWA/y8JVL04+nnuatbCRJcdk2hEjWfQiqZ5Id
nupYbkFKry/aDJiqqzmwC2wBWJ9KebRnEYYmIOu9ufflPZy6vQeW+pwwX+kYiPJS
KNEFy3swvMcitucAEXXGLa6gcq48bF/d5ZHhHHBIh+/7kp0ckOCcwsuOmzfki2/z
JsyeoUAZz2yvNvupH/sZfPInavS7kDpVVR8ZZ0cv5RmxBhY65LYCDJwDr7wS4RD4
glQPdjT2+Q/RbL8Dy/4z8PsPOUecrBXxGfe4hV9pOVs1+3V/TCkyLjNudxroLUrs
AoRuBlvzaWTXD/ohMKO5+rRaMClpLFqC1ADf5CuRxkKwTKYRKUGZ9FYRprKoi9TX
CJH71aOoa8ZYPiPJShcfpTEFhyYqhVyeyapDlyAQ9879mLTLRyku/G9oCSmLflOT
onhMrX6aZTEI24hqHXkU8HHTm5MQquQgLrNdf4iPZyIiKMz+sR++1DI0EWvYt/OT
VgqnPocHWVHr5hmTTL7y9ot8VA0nkJTct9M7rdF7ZG2yAQOYstvPbbf+0JfGRQGh
pyqUOyMNmr48+pYooTO/gS88E1iZA4OSr+Y53K0OpBAH+PXSRlH+KSaAbkBogJdc
0KoD35mFw55YkhhjHkm+B6vvQbmG5BAE9BnaYup5E7Pqz3DbddOdpw6hKZOadqTw
nQ6zp0mY/80AA7PSgFwEAUBemYyGdwpP/B9wOQUol57FC8uz/PpdjBN3nMPC+9ee
aI1xLrVqDDDyHQjKqyj9aZw3ZtDKVIJFThDXPiLSewdQEjtMPq0E32eV2ulvPQDv
wVATtqsyDdn3W6lf4cNQe8ocKcZFUI4slUx0hMzBzknWYrnC//onSYqDE4LDbMEK
KQmMqIjd8kc4YcdWxhbVcCR4Kyc+JQihLmh/b84S8rdWSH5XTsIKM7Zmbl/lZxaJ
fQyLjG1OvW5k/j+BPKdtvibfKR5Q9YEEHjQENAe1dSuwLLvB48VAkRkarWMD9J48
ypWSS/lYaK+DNdNh077lsSRruGpTFDwSBU6Efze4cjeDVKTT0942ugkuw89CFusy
LP23Maa8X82/n0tdoYx/lAOTQ80ftWOltJooLNjvrhAM3RHzAhwG3/UADkuqRpw1
93z5DHk8WlW59CempodPS2geJQHchlMDRdsiIH77Y3gbacuuv01b1AxFmK2ojYJ2
sI0Trk/F7+XFYQD4WPYDOOZ9t9/pgNCqtwpyzg6/KeYnFnrEQ0vcGPnb+w0CQx8t
Xr5Bvjuv/ADvvJjYTZaJcsYG8dsmMLM1EsYz+/cqoAfJ2+Soia37kbg/lUJY0+we
WNb4PFOL3ncHpcxs2Fn8xreYnGKVaC1KoNz5Vksm8pJlN6tJXOzTo/jy3FKosmSy
1ABe+u+RGpqj0iNb7mWVQL02VqMiaBCfiI0vShzldMXEyHH8XOP+osILiqMH9uRc
Yc2l4tHpNamJxlhvvfJqlW+llhbS0hzSl47m4OYzDwlk7myCaZNseeox3b5sWP8B
CJrIxXpHcDtYs9bJpHMVQkArpr3pcMSHq/npJMBrWiVMpKVvUdnwvkIE5DiWoicJ
Xw3beYTcsoUJTQvUF/AmoY++hQ5vYynVtwBgnPD+Rdlqm/p0Fk95gVbj3yR1ctgs
mIbiHm3PoaYik/m9rT4mnhCZqMn4QPV3u2FE2iWr/Sd+P9WkXA8aj+Qqtcnr6zgj
W0/i1i8qnsGhdSlGYL2Vtff3TlM9xymRbI3EjFeJZo3ujMiWF9MqQfR8C6JC3HWK
6ZqAmHH0ATxA1Z+m34nnDxSWLqs3TEXY7hg5J6c8juE6KAWh2lWtZflH1rDCJ6oC
aVpBrIDtBbbqSakeZv7tAl7WH69+SxStaNr0yQSo1i8Zz1DeY1AFx8/SzSbULPQD
C+C//HSVh7lZTLDuv6vwyo8PO909CrF4POX5gd8zJOw3moWHxTlb7CmCFv+J5agf
ccPvV0AvKVOxy8m0ubksouSdEuxUNLApv6fugOkUKmE7BNmgDIJvQdwpYBTgQ2H1
UVvWRnjg9e/gnkjOpPe+FM1VuCZeg/Xyx4F6jd8iWgTpG+rQgRiC1dtocUJrvV0V
WFDQU2jGNi1F8F1peiEiMHBnm0AwptWuF6Ok4Fpg4eL0OwPlKi11cO9DWifWAtwE
4cKRa/OXHbX21QK1SXsv0QcMPr6lMJmfC08Kc2p2ibCQGuYaqvwHfZdtpLBd1/Qo
0wdSy6eubI09K5KMbRtrEdgC8VQF9CSOYjpZ+Tf2F2H0wHTdGpRzwkIhiexACBLe
4HeoylkjI+6TS3SGz6IAyESsh3i6ZiaZ1/TyEOCnp9egtZWPwqQp77GpD55PwsA1
IuSPZobqsCuVTXlXmGps8jdSNqwKGL5+lB9fDqptif1JoKqqV/8VY1iBPquJl3uZ
pntTsOyHJFifa+arDyt7rtxDmyrYbDnkwXEm5VrJTPoBiAygJdESfYrq29Je1MJv
SLoulF1qv7NUM8YLYG52uJcq1iLIYPpDD1VnkYAUhkVwk1Sza1AUZosbsgGc6EPh
x215uS03SJYdbeNAreugemyeCQxWRsdrT/eJDkOb1yDRaJR24/KYOMhG3Mkwzj+F
YCGKagITb99Y8u/qtybtqcoIMyaRozMAM8LvPu9K7hyIqvZba2GAG35inUHjyFh7
Ct17reBhgLcFVOLr4T96cmHLTuUXNz5PJifcSVxBgLmCu13kyJG+t/O9ZGNViBsj
8GVHQzYo3UCqKPW+oFFuciRXWxczdWU/vpYIpIP5dg5MCOLeoG2PkbvItRLPmC+T
Y6UnymQaNKr0KzVWExqjYPewTIkWrhluwT1SaAkIRZ5DHEwEAcEmJrniX9OkIWqC
LILgfTQwklAaPxCFoUlkfhYSfonoWxREePZ4Kb2qJksFnR9BMiRkcQTHSFfadVe+
LJpcgOgCk1voOJQyni1liHg5Et0wvgkp/IJYbSr0iJVVFbo361QoyTL1wrMaEDRh
KQRxyvAuMWWbemTLi/niKrOdLu40QlIXYQHErw53MpBAaI7jxwnfOp3N+4Ym5W3P
UZVB9pEHUaAA2FI7pipy+rizV0xBQDPIBOcvfN6XpwN/VU4MiysjGcgImcOclyr1
VvXbbc4pSkj/7T5t8GMD06FTQO/7wH+R9g7YiWjv0/cANYzKyyAu3DvHKhadzFYL
q8kpRLpYLy48ohbx3PMbHTPcLoLAp1c+7EKRpZSD4YnG28cxIGauvK6D2sM5kcKr
O6ugLiOsqGEJm7R9/SNm/nttA61fdwEvEUbUTT2IAH564LOLLInitEkPPXQEmmLJ
hU9mZclmZPggLW6W53Ogtnfb2rDtj0rZu+0hqK2YAOCHEEAfnPGYBDVxvpPlLYjp
SKbYhi2ievsQPAHZyRq0UNkI31i0MrWByreRS01oD+erlONutZWQD/6oYLFT4SvA
ly+ku0uscgPH4P3ILp3nIQkero8wK3aPfr2WmgaU3O7C4h7LOfjsxqe+m+QJMb9N
7JcqW6MjMsFOSpHngbxYZZB06NyN39P8Fj8QPqpziaPoAiPl0KHn/cqykRTU0se/
KfML5c0iEuk/VVSt8VIGFZqk3pEdbnoxZ5MsBwX4DEdBNKIElzm/PMGkEz+KahwK
F7H1K1N3NpyeJedlLnYgynRwb38NjcBihcrFyIJJWlCmc9LNT3yY+os6fFm5QeV8
XpbMM70atUKuKpANOSsZQU+/DpCd5uEK/5HgtwC059pv/piwtkX7pRNdxXhSH6Td
806b5bKp+W+pKK/Reqxp47fbeAl522wcBl8WpLQK32/Lh37QYxvlMHe/A3x7YClP
ct/7e+DcpxfRoRz6/nTGjTKgRlUQ6UB4Q3+DNWARpp88DDCMhePUP+YoPAKPsTnJ
q1j7vAbzTuUIyKofyQunjAWp+rvOeSjkAVfJpnnDPMeRnVD+bYTVLWYzQ0WAVaNQ
HH9JKgH3Mnwh+T3y2+vyyn53nfdT4U6vxsw4nndhONFoQ/HNusfTFZOGWksz4+kh
HKBMGbjwb0N3F6wPhS+ZLa8FF+kXZoORYoz1B0ipe2tVBx1OEaeXY1xj/Uu7u380
MogyDIl4uPDI7FWFI4jzV9May5MwSIjku7ACoz+pnSGE1wz/lJUSLSA9tYe/Vgq9
9Sr7rxVlG+4cHiMCZLjzgJBOLzgz9Z2zwTlxqwMTNZf1sg/XOeIH/8ix4xrIFlZ/
1TGhWSWZspabhvnesk6LpkLQ8bu6UUu1+jXhO0xbErM6ynnevl4L8DXXbKTZwp3B
qhHUPnvA3VNXncAQ/+bXQ85OfiBwuikzrZLyBMTSMREK6//IvjgYqamVmS3o3Aj7
6+2dbrf4lQoLDjHtUYM9EWLuYSZJZ1OfEp7TZptu9sIiWQH2+tsgxiI+l+bZEwM0
XCgD/T2Fc13F04bcWWFhfq50UjdGfRu2p6cT7hNW1c2Az81fJpeiQ5ofOoYzI17Y
OQJEUSLsvyj7JWISafHPIzjl49vjYjQ1oaPTXra+YiEs4HD6SdQobWkROyhcm2L1
uVGp3MyN6xcHXbhrcK85vJrwPNZRVB4zMVsw5ysQp4dSk64uvWJMvfwLtfTV6Mjx
Fft9CIhX38oOP+llPkaFkWnexXWpn8Nd5HnqHjuv28x0OLIQ7LwlR4QXxOkHKlEG
14FTfBSKu1of6W0HJ4UtnJU2J3ynYDJfQbGuKxE6xXjXKHHNVeZ1Q7sg0URR0ezF
VYJWcobowjkahXB0RRa4mzy+1qSkGQwiQQCf+bJfDFtDVV3+KKWC4txgV8XDsTC6
c/3hyl9Sedmy1Zlacip3eQIlpJn1uqjRQPdKMAamrskWj6Cd6Mgjz29DOZCEDBCy
OQ8dx/ruiCrlFb+xzpgHrrT9n/BxwfAZRm0OznSErDIsdXbD6tUfSHf8EnkAKwP8
KiJw+Yo7h7eXsvZJpGBPxzu9tBznkr77bNzVzibcQWN5JEtHruKRqbpJt1HmcHFo
JJqff90VQwMp/6+jS07GqLXc62UfcN9M22h0ReMwranNl47dQzo+TRr0zOoz5Rb4
ltmit99x37I8shOyzud8k3LyoYrZSvZGd0jOO0NNXs600IimLsLmasdW6h+580fP
W7ZUzUzjb6JVDlYFKS+xUjLpMJICiLIh1ajfvBhM7tobXOR6/ZcU/bgFj5eD1hKR
jSI6GMJaXN+Cfl7assiQ4B/E2ZScsZ0htMtqDx0kK1VeTWr3oSzFbh/6r26ry6/z
ogGqsedH4QvN9n+e7foDfY5OGkGVxkkm7HW5f9RzS+p4IUF7Ze5i311G6J3s7CfU
IQnNcBQZVx2WNxjg+Y++KXJiiS2di0hrLOnH3vlI/bBRYmWchiCCriuAG0B7QqVN
PmkdaN3FdptGBo3Ou18UAWESjYxEzujRExh5W0NpOG5CIUaU3IaU90tYXGtCdjw4
45wd28xRRSd8x7ZfDrVie4mXE3F6A1/M8q8jIe/1Bj0/FwlVtp//RcUCap1VlQZU
XrUslbMMwBB2p24VNJGMrBbnYDuy62UipXE0PWo9icFvzrMJne+d1u9fzwCKXC+Y
7P2XjO0TWfKixoxvk7wyfYOO0uhu8Vu76XE0H1bdp0TczXUxY8rwB+m2D9hnBXZl
2Ydci3ic4kgjsLtx3t3JQX11Fy9DuE1+CSD6TOSdysu5jMXX19pptBF91nNKZWAM
LNy8MzRN1paIoFObxTelNISyBjRQzpW0XqPiB0Gm+hiFTwlXZDfOe0JZd5pZkyBR
6z8NdMpkHCA4Om4cFz7wMEPAH5ZWVj7GadZ6RBCJ/zt6JsBbHYjnhK9No1pCgpG1
VfBVirJP5aSYZRo455GZD654aAaoLdNVAHgCX6GC1dCP+KJ9vDN9nwnkrIgo5q6k
PCJP+4RFQckhHC2CjT2qC9vWaB5Rub23ZSW8atzzJkfQhBb2oK92tQZwxScOPqkX
CVOqyesAJDxHYbV+97OVaJESJY3px/odsDxGyFZRJ8a/DSx4AOlQKsjQu87OWAL3
DXEoImtPfcLvXUSUWn0dHAVfhAOtzZ1TEmP7TZiT84R/9ZL4MNs4OOvx8JSkHPzM
WPquNpJMT/1ViBuUbs3yiFx+nyMG+3alkE7qEffDlO4h5G0a7D3xOfhqaNmpgyCm
BDakdVcJN9nKyY/LCWoeq4p8f8AeloiX/QxdhTys279CkB5YFyXvSEriHcaHhbkp
71AQv5D2cVDkSxYKwFsdf9hQJqsrm4x3QGpqZVyz5bT1dcn9AklFCjcabrgvpdrX
5RweMaI0Qz8a2PWqrtHlpv2rav9dw4yz/V1R2nwX0qx28jAJ5BPgaNZiCV7F8LJF
4IVmR4ySSRt4kRBegJqXqoS/qye8s/kjEjpe2mdQ4IwLwvLDJq41h3FbZd76OQbd
Saarvd/SSchsq+bqvIOHfUqNbdiBYMQbBIXKhL7jdrBD9R5hsVVHFau0nD8YSOc0
gGtadA3talOaUlkQ7e9Wjar5PunBZ9PRE24jQE3MIW3TEu30SMSR+K9wSkf9FgwQ
ZFOpIfGG8X/47ZXHkixFySwrEi+O4RqxaCG++pB7No6mGYHSzSRXP69h+I4z6KtL
+3nFlLNYbjeT4s/t0KfGJN8LuxRyo15Sm6HjYqNhCcJe5yrRq75x1+NfPrWwqrAg
uOg5Lc7jC1tqEYvakJnOpqGXT+oq8kkbO5NY4P61TncTkXXVYTnSTBXfhWmfhinT
ujOB+rYUhEPaLOC4VnQgO7jfNrMEyaMs8imkMnH3UTDjmqldC3KQuqf9WobZz9rS
p2GFch47qxXhPUeCgRBcTSjkBuV5v9/ce/D3298xhJBzF7/YbbxZIhJFQGBsLvy8
t2BSmfuBo6Evvr4ZgKebnlkzOcG6FGxJFaupxqiASIlsf1OiNhxnjiJaP1flvxci
CHzNNYBTJa9n5HnoeJk6+n5HpRhdGyOZ4DpoNog52fkU4sMb0AkkbNLNPWaOx35Z
o05qipZvYTVPdK2MA8x/SJTXCs48GAUzYKAicetdpDAintMt+CS536y3Cck95WnK
pSmE1nZkKSvm6RhE8axZxDCoPaV0f4OnOPtH0ovpJvZzSHgdNThZKR5mo2Frbqqk
ove0ZMIYk43Q1v3INkprZE2LJvOH8GOrhbDqB1SXdmw/m5brtT4e1UqksUIEtTPx
xs4yXNcnT2emkWSKYz0eg8CvCA+idVYKVU8OcEXGiHBAfa8nyGbK9biXpiRKR44I
AWcNvpuuuTlOuSmLV6b4t5GZw+eOuvCBj2aXn93AIUw+edhNMmu/61Q/KUmB7EJ+
UyjtgwdNPRzouYMUxrcoGs+AOiNFRZsUvf/utGXwt6omilCuacJ5NRU21xsMdFzf
6gbFuzl218FTzYH4jqxuPHJSRXy9HqEvHjhL914mDAwoGMfmZB7Rli5EQHwiIuFi
fa1eiS0S4aPnGL/ZaBBmvOENJe6FZyzv03I9hFGlvy5R24Bm23a4NZFnzQ1IPT/t
i7P4crY570XsLO15Ffpo0tF3h4lSOerH6B8332IFegh4c7ZqK+z7tmdyWRHErV5G
1ODR9g5NcRy3R9+yhvHRm5lWQntpLaXsD3zt7zsKgHqrTBmPPKOsVMzWNhLC6t2I
sfL26UDZ5ZonwQNsT/3J/9fulRA3pPp/7qMhz5gGQwM8mn/RUwXGwqGqpaSO1DYQ
E3Aw+GP73FaE46rALz8zwJdkD+wULDIKwMQEF0B1g0CezdHb+/OiojHmKreit72Y
LJKLn7ain3U5zlHmdIystrFcnNpS9NiIpDMftKHX0rlFNWV0ZnV3ZHVODVF6hjZP
zJTwEyWMulRgxkuI6rJ0SzMQbWbY3xU/yh6doI0vpS+yWq8U2PfszpQMRfdtK9G3
RQ6ba1hXZzn2IRNeabQCFs940D8qu+3ekkCEZSVLl5dpgLCSBqGQLkHL9T+jq2Ua
Xc6aQ22gwJTBP6zUeQDKT2RPZ7ak3J1MTYeBbMrFc1HGWIppXgPa2xjzHXuFqjuy
iyxuQUOr2miTIlmgpTg/o0I8RFADFNuNFg/+6KA2wo8/W+MUm0Nq4bw7rNg6XQnS
2TauKJFC8f+9+p/2saoTSoGbqtb5YQ1KHZ3k6rLVsQIhiL+8jx2xoU3Ea1M6WqIb
B9T/Y5iaO0DCNLp66O+DoiET8C7zaVdeHXUSfSgpM4U/Oyw5i7hc4QAZfZGmQog1
73tGiJVE36N6FDhffLBvvohe8C6CZ2V1oXK4uh06PLwA8uAUOsAGxvKSU+YcHcek
w84XflACTWkHI3d06QZO5oVPO+PUHK3R0GSWKoWzjPJij9C7aBSE+eIQqd8zyYHB
F6enXYQO7iQ0RZvk+fJiTRw7NgRGywCQs+AL4ITP+aGuD5OI1NnVE3LBuRbHIwWi
sIMptnptbn5xQZJUs5UUkXL0JFhNHaB3kuQVvOkqiYqK/Sc0HASYg22RDbo3WeYm
0T3HVTt1DQogoeu9EeHhuhbMHGtJPVN4AeGN+dnpqi+ZSxdWt4h7DGTbPqMOVp6w
ahs/cQAhIWon0gUuAimnOBgVK333lvjpgy6EUeYpY4/7b7eT1Agq7mVI2yD+g7Rd
G8d25HCP20ZmG5dnTxztiRVchedghlyKpGY/Z5pwPN4Ooka+CJgfH6tmel1LRBPD
UwzFENiE5mSCeT0h7/vilXidUIHBlTSEQEqTIkJ85CCrUrRtqF3wmNylWkpmFq3j
Jxqs3ogOx/BKTjNnA5JpYi+Zmsez6Py0fW5WpxzcUxgZLbHLYip4sP8oK3UP05ZV
NAtTeNk7Y4q2CsxM75N+bEkAE5g7AhFbu8is/i0v1mEthPSsnN5kUDtUtER+mR8Y
TW25HK0hxsNbP2tpn4k7xjMlFOnBuZYX8J5ABmiGsu0oDSx8PWfqU5eKNiT2Xcp+
j2aqOAaSVLKS7OcLbLw6LQZTOdQpFfmQn1RLSIHvw8VduDIxoUSUFwRtmqnG7KRC
Dure36euEhoMlNfr1BSE4/sJ3dc+S9SGZuAmEaLstPAcacesUnrdU1cUQYp5eIrY
WUjDUqfBqI4yB3QYzr5iQsetgzwFYL8c0K/+mdNObo8JJ9RZDfhK2lEGtX7MNHpB
J+KZ+WUzyAQl5tEjkzU5hYnBOT/WyU+0wibaaEqLgoNMYmLldDiFm4Zbk2nTyRIo
8B5iyE9rNdlVef2Vu47yO6i7OfH3sWZWlob+J5kxYhaxcS9QaYJyNhl3gATAWWVb
dG0a67NS/xxHbDUVJHBAnLL2N+xOhzEh6zPczVHUoKEnGF84Shtpil/eUGDdlhil
i0OT1cESiBIhP5CNvztJ0WLTV9/E9Ak8saRfmSlI/4wp0xgz1z2tzz8Q3SkxKAPn
lL9zXDT76xjDJzwJu87tYtdLkBLBZ/Iu8KeZfyAcKBeZIiI+htrEIMqqyjEH8OQ4
b8dWB9hAbGEnePbVTORS4Ajn93J19kXwY6LpUlvM6ox5l5QbJoWLMgcl/dIC2Sq3
vUz5e0uEh93cl6Hjk9qq1eDKOu+z1SEk9bmbdFUt3AM1B2vt95Sn8CGOPJifS+9N
uIVSDM7IMwiEtloNjGYLYWufagXaLw/GntG1PkPaBUtgkEgaDaD4Fj8ZKBYvDJgZ
m3frKEqGzSef6JFq3WiRqn4of2yMkIeiYyxLj9zlIWLZt7+fvIzrlV9eYo+Fxdlo
4caDcwen7+GgIafskmr0yu27A/V+2knToMqbwWoi2+4BJrgNtyPRZqYZJDmOza9i
bUJIPKxTecUozSiTmWtMi1XuTBR32Pq1vsfrq4iUk0J0pNFcwWpK/uohOA6XiR1t
2hFqXrfnyb3SqXUxHvQfLWKuKyLfrxjWMx7Wg8UtH6i+YO5XP6mLKAwccLkdEA5u
mZUyLLtx9VDlAyXBiCY0zMQkWV3uXKDp4WQcUFQPgSAU3h4DkU1ANXNWJYpwGe4a
SnGKgVtMw7k9hgakgXTmrWJ+XwKih2VSkvSuqAHK+9Tpo4t0y9vPZHy6rSNc/xY/
BCg2dArHsu8GKq6zs7rdAZ+QNnqioEn6FcnUvjPTFgW2nGZKicmJ0IJ12rWG6/Li
brNzmB0aNNGzm4DWxNlmfCc9S9joNWp5SIgRsqc0GVJQD7Av55bhG8E5eUXpKRPL
7MfESt+UBB2kdBljTeATM+XH7QCIB37ZgsXZecTKLejcBdF6P+EetWoFWxVZQre5
GG0vB+x4AHpw4Rs10r3IrwNRBBjXCWPrR8AwaP0jZ9Wpt2yveM4mqG0j2gNLqOXJ
jWCZM8ibJXtFyRKeSciE0y8ORoVdEFa4T3IrSuoA/mCeO/4BiUA1cZSSu4K1Hm0h
lMYIAgzWRI4sXtIIclhjTkBKzq4le62nwCjirLQeUPuO1LR5J3LNlhOR7vaXMAes
08u7C78Le5B3BHmPLvdWyapXBdORh5PVz6n5KrvT1UJHJzNBO77ka+FSZ/qw4lGh
uVYC7Am8f872I1JCSe9KDMmzJjNai4IQ04cPrnjcDA6nLLxLVSCex9mpmaMMLik2
iqY1umFOMNvndy9wTcgZjaSXDfCMwuWWk2suszs6xX19oMFLrtBAMbicHOxpAVio
eGRBbZUZ9vgshLIKPsZb31IBp/RoqPIvHpaUxBIVWoYhPisYNHkU8JcHEwUuMHCK
JccCYOlDPulxoZEeRDsTUkYDy62WHC6KpTcLyQhqbjhHRN0PEQhnzKyEuVwvO5iH
OelUZJ1EQQ0aydS6BBVFfvnUIHl3ydIX5FoXU6DEfWGzI4ujwwP1W6HCHnIQ+lmj
IBuRmSXOGVbMROX/vQ5wQr7Ti7aM/BVqChRpqLtgEoI8MoAPkPEwFXusJoNwNnFp
jGuIbvN8RengsUzh6StsAk1akDjQXlWLhNyfqJaPQ6DN2HkheGqDej1pX2zTs1Oj
FWOOkUFj9lOpNVcWbPu8ECBUJONoDNR+9t9VOrc0LFVFfsKL1kdy58/+JdCZOrEL
V5H+JRGGAWPTPMd/ZHcHzFx0md1S4fqkYLEe08AEmCTCr/DmZqi0OBYr3zLrTMpA
4KC9UJsyjbuFsaxrRo+PJV4L7DhMVWf1oZ29JtaTAaVpQqdUIqASGkFTFWMD3N+G
X95UaG6qBjzVVRWz27QMUn8C3Kv6CkUvJP5vZNONmjYwcNqng/f/wEHMI6PV+58k
ipd6xXndDryk/qoqZQIXHjTGXyNuLvuZgcLRGhabCyqNOKp8Mzb+k+bDKEBbzuO2
jy8wXDeWgdekIBljlXm9cKCdXJdMml5aNLyVkV1sMHqXN+hicwRBRys2gPfUJbMW
cAWjigSazxgoacAFWO3TvGTqEVrfFHqryJNUIDX7dVcw+BZ/YHEarV2u8cxNkt+h
ZR/Nmt9BPs0IJy1aJMf9e1nU9DhvB9Fh/ZidvoJbs51dZmIR2kBXcE9WLawPhJ02
M/LLHe4V/GF9aHfv84QAqRjvxSCkM4tlQgbN20XVRPQYPi3M7nfLMpIhbiZwMAcf
qAMFbOfbftdY/Y1VpLWLU+ifFAxPnN4W35IALw3GzuS3JEJb/3HEGpqodyeEBpsN
b5CGyypk5AI1Aia9K+Ev5rYmNYMWKPHeYiAhYaQ2RdiJ7P7cUxUe+8EXvweM/BGT
Dd2QcvRyGsqsxEUskXdYL4GMBj72kxP9Sb0l+LpKyZOgJ4uNi/OHOPMfjUSbnlho
MBHvL6fI0AASNYj52nDnlIMfzODNy7fhdspJ/RWrWPsCtD/agh3hoo0qNPve8wkH
+I6efVbkLJ1SSYNznmHJXabQdh8BUNMcl+53F8hlxoZ4c6zkmqI73RzAP3Td0Ukv
nikEAqE/dNOUBqEkkPVl8YzyfPZOwwJQjftSPBrE8UaBF7V78GCrzq5IquoZ2aA2
AAP7m6UnAfKFgHAkr7JpQJ8lE/zF1p2uz0o2vXoJei39ErVz5qhe/vJYsI3n38QH
CKd7SY3taJkuDO9hWTMbMWptFZxWclsdz/oQ/FSxEyAGt8GRB5h/0Ldu0+Ov0o0W
dXV5nL8hfQkSzTPdnuOztjCYltui/iBKLC5oYc/mYzfTklyHtUEy0KQLHD3uTqwX
mcL2XA/WMLsojhLZooXsLLl6sFk3FBhDMOeQrSTb9DrFzD0sMl6GNV8wKO5EMbK3
Ym3Vt6P7/kjiT7ABr+58joYRsdzEIkIqD9boubQakn1lkIOrdkeOLcO13pZkWTL0
pLbqzHoNRNFqYF3Ah/GP89iKdsyFsn4BQNQ7w12TAKpNlL3Ur8qlIayni/+6VDc7
6G9VnKxwqLG9xpG2W5zrOE5biGq6ZAjo2/mlsJcsO6olFi3atVvmJYdpDAKcKhFT
pX6UuJdWBoFEnt68PN5A7pl5Ms8LYO2NMbPah5O4G9Iet8dGupns83YCPUR6ZkaY
vW5Gt31POszQjaEzJXJHtg4H37IB2R9iLrqjJv8akq7qZqNCsLF0YyO9Kl02ei86
MPpsAQt+G+uJVos3zRt/zHBhsApA/QTfn9a/8dIbkuLeqM2XzOdKC5+7R3Nxl9F5
zVNjB3zoU76ozazqoARAGwUsR3vG3iDCfVrcGuplm4RYDkeXnx03b68rq8M0i9lx
cTMtH5XFE5yaz4bbe3yENzYjfLsPkpHe+slAa03azLu6P1ZL9U9EW8y2Mpt3Oa5h
4Aeiz7RgaqqRUKkPhya9fxQ46/xB/mXN4wtKK6DLUeGNaIUcKpgYDIeQ4zLK6iQI
zqZndahm2NlHcIiIS+dBRGqLnYVudpVnjh8ycl05uYrnVKg5B6OiUZDpe69XU1Ds
A/MIEIO6i/sD3ON1kLVC2L2bjCjPJEx7MMc+76S5wSGIhORiHLVD24nzz7pct5+f
nKAuVwjvXpTBcOIpQs9/PaS5T0b5pL9wz5pENz/Qfboyh/GSidgFBxHOr0syBDZB
tAA8sMA12MYWTTGnQm8Sa/nAXJH5cLS6CDz0UQXHiTsRbT8CUUV4QTCgYHRyqiGM
iFIFxl+WYi6oZ5fiaWfh08fax6uu2dHx4/Zs1rRGgxE7bZtikmmo+iGdke4rl92M
Unmxp7hRpBx4TR8PTn8+T07Rpda+6EMnpdLGXjm9cMK5eAi3rfWECCt34Uhrm/tw
chknh9r8oL0O3odEfX8+hSK4BDM6n8iBReIy09e1p3WDuiaaGwDZqhsxiaGWc7Cm
CQeDir6yux/emGiwP4QUExixObvfhOq0DH72SaNO2L7RAQw6yT1yHAG+9yPuWxNB
5Tr8oOmhZ7LZB5Yw0YC4sk0A4hVSpzwmpadgN+8CJ6itqz3vaC/uTDyIj+gWvKo0
Tdu82NXBerYApdfPDW0/Hiz93/J541/owwEiiz/K7KKH93nb3BUiOhhWS5eoEfAw
KiYgSd9OWh4AhWSO2ykajPHEB01Hi8OXKRb5foy+l2LsoK3heLcByQGYa5vMiR2S
ZMVdFCuQFHjiJ1Ws95x6hRTapDDNLhtUJbf4yPhsdL+X88awEYTl8zylhtHpmEq6
3cPqk+dair1f1dBFRSlMOM2l8ktFB5HUsDtRCk7kTTQoSi/GEgDJ7XJRMAWraImc
akw+ef9ksdpkrE+5gfV3OPr6yfoScv/6J56/hJTcCcKRKErWrOwHqhn6IGeuq821
E4PeutFfyfpRM1hT7EeBD189Wnt1SYsSpTRS3pH0SIGhSjx+gsvt5tRzTG9Q8EDb
P6VVyMsupgLsJuQ3yWjdJVB1gdVowf21BHYMTHho9wOYjqgHuuOVu86XEA0rXKYE
TyNfwhfDm8TmqdoSFT25PlglXdUbukwSJ3Eub4b/hD8GIZNxkt2hvsUySGNvxFLC
YszF9A/WXP9ypcucPpsj1sG/x8kroMIf47W6qtW21SSq77WK5yptAttng7j3OY0z
0q9GkD7HpU9aR5qyMKCcsrx9nnmsDDIuSTJy6QCA1UqDVXftB8ypuztz46nyoZvq
yepzG5+rnJ+QmTd7FvatexPfga2Si7uR9lpZJP63tpa459orGEwW6aoIuOT0kxxm
z9tJJf5wXuCZr9xbQF6FW3PmWCksgGvVcKOtaHRkht938VgPDhHX1MHNp44vJMDZ
Jemsz5ZqSzGxx8C2vPg6Oj0LSSWaNlGNlOIlr+VKm1wGvRRUz9u4zmZNJaz4TdEX
NmDf850BGItv8liE11bim6wcVMiO44neGk9j2dGQckxS+IuJvIgf6q1jY1c4dPY2
oDKU8aRUDl9nnjV5/MG44rI76ZeWbD5ty2kQuog2WUKUnTlXW0ujkqPU81p62k1F
2kWF/b8vEzxj9YKr+Txyg6bkur64tkxnqBSzhdYXiD2TUMcDNCmdv2AoEPHLLzDG
5x7+TZ4+o2xhs1iDY3Ri2EBfcXfCmPUVWZVqKn2LCbPDrTE1k6nht0ANGTK9/yNc
QZbOBoMYszPkMqtQOzftvuXkL7VL0dlEl8jxNmv1G4gNufoFyiHmMfcb6D3A+LQf
1fqzno5iTSC5q04ZYZR5lBL52ivyW/GJ2Qq+l9opTJieA5TwK36+beoJ47LCVx7O
9tm//UjvNigfsn4UPis8hcyABFXk526Z6DsJNuhNqSRKFm4xodZmtavo7XoeLSC0
eml3Y0lxJWEMctAzKykeJc1pXZOzNEG7PuQggKsz5T0fPVN/LkotGkP0sheOrct9
aX/ComALVsK2Zoa3VTlzh0eNa2534Ysq1VJxeX9nV7sBozYqiKrCPf+dPmP61bPq
2ecynHffNT7CydlfJ/Xxwj8zu+FDq5RanvSoRqplAfENenDpjzHX+1GjkNoXq6Gm
Mu6ZejvIf6mAJS821XC6EqfNMDyQtTXngBXrOPSjbH2/Ioxrrer3bSWSdzRLMvkt
z7C+FXfM7jefwwJMIG7VQoQL+Lxo8f87RiyN4L1A7G6gk3M1QiPHDZPhJ8mo7bsG
yZKxsnXJ5d89M0MOmCzYcV5AX2dGFVEoQmL8Cxs+qMffqNQT3M5Z+jV2Dl8397bM
uFAq7r3nb6NiDIjXDMvssCPrvASplg0h7KN1WOUtk6trvXgle0FBF6u2rCfdwie2
AO4zTBBry1zXg/dhbxMMfrfNwKPXUBv7lRfM78eSIq9fyTW6xCPVPqgmmj0bjUXx
3i52bdifsCsHdUZrMtfygQV/TYKJURHOpLgEunjlGwKy6O4K84N91v+WqafKcy49
AduwL2bkQb69eJxFEpi5p9/i9tK73+wywyBSMfSZj0yOXMQaRP/X0ORnrd/GNXDP
KhKiMtEkv8hgX/axVSPIsnZruZP9uLWwqUz8DCGTG+qsjA9HwWULwM7wmEibtOrD
AJYRJBYogzqoj5tJEJ7BUnhoBhxHqclXpxXeEZ+/2/TfBKJhEFgAjZpVmDXQU/jH
HMsljr4W0ayxlNeubNN836B1GNbCUnXGNygNYdMjhrH7FeRk2lMEEJiimfJrT9FK
q8vCzcP2EQKAVoAxCP6sYu9ak9jRHFxgy6bTtMEgTxAcfNbEgLBv1r1D5y3zlw9w
P48xEnJpUZWFAzNvhd8wgBqtkBD9+6JdWHoDvI1ZhUW8qBUFQkbfWNvPX/aZeK8d
50vVx3ox8Flu44Jqo2xGNCVpNfQ2N8MNSfSPR31bfGCFiE8kjX2vnZYmFRKrUPXy
p7koKOEoT9LczY8EsYz00MGdXzXyy9xgiZtYRcfIagE76Qnd7lHf1U8KfZlXrzvA
yaRD5sGkcE4VX5bdugsbAr9iK3WCHdu5xym3oczThThrMoyEmnZNt1IeO5GBHdPB
9+7/AFJqzKvLuv/o/X1A5fC87kdrlma+7hjG36lDw3hXrFEYk623V4M551m7t0Au
LngIuL+M3KBDmJlXWAsxCYUfuvXBYmDS5LRq2hTRmaGTiZME0ZQ8mQzgPKnpEFtO
/hrSoygY0xYTIOEE9o1VXDcs8aivAnY0MIfENkUNnDVvA1iHKy+FQTleI9AkvtRq
Gdyke4+d4ZlQf9JlV/t3PYreXyIaU/U+jgBvXukPkRlkO/r6y5gD5Bje7Xo8AWAx
DdfUFo26phoG+BXrpUc0wOGbBuOY2cy9XTW0pN9v6sY+1cQ8kWtr4WPo+QgWGsnX
gx+CxeF0EWqcwyNN/u1ycqkXdJHyKnel6WCGkcp1RuL25jAtoxiQE76TRzUtZd7x
tQWucZAen1IVX9Y66fVHjjLlnc/HDebJnqWxmJpY0Df9XGN9aukq/QPELIsCfnNY
h6oSfnYodU+eSB2gsUP2y1MnWDhbix3IuRKw0PgjoAMgIMFfOppq19izK5RJDAnX
dMjcY//gEZWy4wUm5m4m5/lTt7SQSkUUEvjjviX1W1KLh4qoGCh6Y3KVgs7+KHQa
2MQsyg43gxnFWH3z6FDzS+U4YuCPCKyghLXepNmKLmJUb/yfBdkGABvHT4AU1fp9
c8aykD//n6qQFqRRjeuBVIeacHvcjPu2P9KMwTooCcHhnJPU3aYnUTZ7me0xhW5i
mADdKSnQkX3Gjf89x4V9rZM2GDtdMkEK2BRwfgj7IELvOtLXO2JgQSv+mlAY4mS2
Q0h/CNql79OL8PxXjPfaI8LmiVxXgg56HH6pECDkeR33XGEOnYlkrIqf0LPDe/hX
kUm59iN/p4WQDz33Trqj0y061h7ir1K17KabBRlb5elzgGThyGYA6WDTp4gQM8j+
CIx57oSws3KOgFQwNxe/tqaVrRZE/uZkwv76cV8FCN93QLtWGaxvtBWiv+PPP2aT
zGOGkf5e2TnSWw9L+sdssPzojx0aB98J4iW1vbcRU4234B0n5sBw6nlQthAJ3CNs
63Ln4k+DHuQx8xyCTdWU16fRCKBTF3b1lJbAZ8puJtREfihiNEurtnKnx/vsqAnu
wqiZOTMVOxoz2prBmKK5Og4ZsTqNVCTkFtSEDAtdaYPxTXta0MqCJXmDjlOHgQlC
0D2eo6itizYfx5g1AV1DeHoKnAqhZ/RltuPhak5wV81o63Q1u050AUgUvez2H4Ig
bAqONkjHxSItzfXUF1arFFFIfsMBmEK+nEFoHbzjn/CUnawa+iIAd2a4KjWbzRiU
lx6gvj+Edw0UI+f9d/eogi+qJ5EfG5p5FqOBX3XEJw5fi1WrvKI2ml041c4gTtWM
rCDYNWeIkQuKfC0FuTb22ch83Z4j479nYkwyA9tV+Oomnhz62B2eJ+tHr7bLvaj9
SR6x/3G0PZ10zjV/S1da2eFccslX8oxu0nAxGETPwLfp8AqUdeu8P+KLreRHmXQo
Pt01wjuRUtbjtWq0cDa7sVKLN6TiTbBqrfyd0cEeO2fsSgyuqf72aN9I9mpHJieq
phyca9fIAQEWsaOMLanexLwKC5OtCxgoClZQz859RcTeMW4amC8xalWC1LqxCDqe
uMm9SQurlaApS39aW0PLBhPY+Rgt3AwJO/aXANAm5ZZ4Obe7+n5XkOpO+xhRdLwx
3NjX8TXOgXSNkB9TWAhTZ6u8rtNGkqaKF/mWs8VDTYkUwbDblEoDqRXCZPh8Zvka
xNInUmdn9hHNXWFfsqij8AREebt0Lek7jNNfhjTnwQZRYdFF9fDXAGKCRlK70UGn
mWcOe6MSrDsJIZQ7HMM5C/rxifqwNRajOnXT0aj0b9QOkSR2z5+9jwXDwm1+xlEg
4V/Kd0JUoikHOadioR0PRCtH+iDLpBUw6f7dkBvSwDS1mTb7KLRjXEkk+Oyuof41
UtIU/8SzFQpcRcbiaWNMaVvfN2TRTnmw7Tiv9+TcsuvuptlSsL7bp+ljVJzzRza6
Ysffe9N1iRrP6JJr+mC6ebsSeGaoBg8mC/rXvEAocLvy81BeCNv5qTMc3o1hdcGI
KqyM/tLrreO6vC2FECShxNtR8hKvylV8CFdzfymO4rANzOzDjOJwSfj690I72A0m
OGZ3J5Qx336avwZ05SlnbK3bMSmHAKHuwbYc1Bxx5B/Wsbg67BrSgUhm7EXplcHz
bD5Yn0nE8fXKvC76hOX6mdbRbITxtZ6QEWWbkW+EekTSOPqzeZ2vARZASPX26F2S
H5qaTXVel2+D87/h2HT+48No5Dnrc2ViN/vBy5+vSyW36FVvNZ2s7E6l7YCHPinZ
n8zBQhkJE+FIoJ3hF74BYtJupgGEFxTj1lMwaqcBXmBhLCJAPg3pNlK5oidNTGJL
183bEXHWrAVHHu6//cwbRXVI0Nf/4oFYeLEwtJw4sPqH91hDunKAny1RSzeYAfwn
RmD+DLCC2DvoyWGFbsY34SFFrs41405txw4zb7fOXSWPHHTbMIr+KpVatQqTIMXx
UPNbu1vhnYiFylbEvM1kdAYSS+79Y4aSJHw47eIqSxcwco0l20xc4wfOKH83lUte
h164yRIilSTxMJQe79G2mpMFezo1dW6vsKdTJGgTfq6HrxSXVsilyLI7aKaMX2fC
aLNwsOYZXwP46/K3LCBC47dCtE7+Q1cKa/7mKBSF40rgn7rKC1jqwaqoSXmCFFZY
ig0jJfmOfVa4PJYsL3j+O7rPPfprnkefeiZCUBtp/n0vyc6+NoQudAZrf7jdf5D3
nPfOONt7TweRyUJ8IZo6C3yFzuX88QNu/1euQ6rxhH+J6iOjbOxgU9jw7cNbFDeb
lKGD1mTUVpWVX1yu193B9d5bl0wnv9LCX2/Qj3uyNILWdZuIrlCnM0BIeIedSBMA
gmQsf76GZ47ZOMdrzd/gAtueOEIfFeeQLZRGwV4u3zQRluBre6SZJFTL5PmZsKAe
JYVcMOf8cvqbjrblQpz8BYle+QqFZe14LVFQhettcIJD17BfZfTN8XECk5nsylrE
+hR3FQt6r8zIi60ImitC2JloTLu4EGreW4YxMe+GaT54ymWtNTVBSWSoPrGn+Zhd
ujT+bAiSQU/CIyT1UQ6joenqTRml0LRr0/ELA6rrnvozrboxMtvQwtDz/sEgldLE
m3iA8+sERWKQ4zZlawhQh2av9OzYeneVeC/JHx5aEuZqzwAFl1GHTp7QrR9gcSgX
31sTLbODuBvM3ldTAWc9bL5JuYuZmGnDj9eIeuC/oBxeiwfkSNUqFYzBbb1h1sj0
k1+MV9G8KPKlv5Y5HcM2ch6X59eu0PkVSBcAL9KR/utnSXAUiSbGVu3D3pNQakUb
nJ0XP/EUhnIKNbyXiPKR6EZSBIUk6JOqNbWs4QYziMQmiqLeSVMTUvMeDX8eNOI2
HN0ZhlTxfJm2bJzXZcOSjUAfiBSTplrrcON2UQguxCcMJK3WJuiqbvY8qs8hkGI+
UymEJhHVt6RhQN/0n405Y/a5yds4bjyxvCXJyIMpp2IJT+D06EPxuCpOOl1el/K1
QPlSw5QZdRkAPV8lzMPz6RX8k4AS0UEtaXsOhZxb4hbnlUe3oO74Jwt1HA198HeH
IkwUVLkTvjSuJ8UhaNOtOsMDD4i9VhaB3TOAM6ZMUGQrhG2puWH15rvBMpha9pJt
H3VRd5PkNoS+1ksUXGrP7DdP1eubcG78Ljm6YC7TlmI85eiqjg1acHkHNUbRw/Na
JLwVIVRPlAfbDR5E6QVsLPeQ+mCvrfFEItA1314GXncoStfsEgLeTS2+MPZt9xNi
yYu6xqbFNi7NgenR5fPz4jRKeGHuEpAelJSslCELBFslSUVbwSmXmrRC2ry3jWvJ
h1qoHnQZR4ENqO7UJeClaqxNlJYDeDjtPhomSMV5EUV6Pp4fK2otTS9fcKJLzvSw
gHYSKl/MbX4+AeTaaE9hAtE03GKsw3CEfYTFHnYKUE+kxlVU1JVkWZ/5PEtia5gl
Jr23PXPChHqRUKpcc/joAuIMuIPRCpT6iCy8P9pmITv82qF/Uy0NozXUCZ2nIzAU
GdD405LEqrsm4lbkIvns4a58EaMkECKe8FidCft/6cCZoMUaINU6+bWIjjHe/C8l
WNEmaaqPI7OVtBdcwZhUlIWMOF8iqKAtKd/HHgHnsv6McSpH7Y+W7e/bhGhekBb0
2u+cn0ptTFbmZucn+d5OgIlN6W93JeUjWsNZxMvFgde12stSjt825IIXQ5IVn41y
daMVngs+OVhptrCJTMIBzvoSGFtFlYKNJEjl52UT64NFDUiKY8r72I9ZeN3kyiTK
R2vZZuYu+ovQULsR5X0MLsQtdkFWb4bJhIBzpd/moDCneJSGQF/gRDJxG7NHCFk9
Yoe7VJJrl7x+pH8xDn9Z+4l0JfNxhzssOj5LvndR4HRd0Wr7ldvle0ptr6gUa3SB
PYFfqneU8H8KZ6yl3VLF3doqEXe70WrPiG+UfO2BgOEevV9ZwYe5r3zMkToVEqdq
Xjukv4CfrbDEOgn+nAnTXw7k0a8HWlhBxTwkr/M00wBxxnSpAclL15uuEDXEsXSY
SfmJjPr0hHORcXY/q4cqc1x6t0n3pHYY8EVlk8Bzs7zAbMxQvtPSjkksG8pAQeXm
0udvoMcmTPCBPVWDMqzL4iC7YU4mtazObS7bbxebw8xF4mWhyBs/AWU1Oh6dJbp0
3lRJbk98dmNizomDvebGo72NPhzxOPJ3wbdoLilf7qtlNdVEZtzGh8mqEBqn5a//
GU4sX7Lg0tpao9+Y/OANYDT5Xts0cPP7zFnmWTuO5NbbjdaAtDyUcvD44BE7d8cn
31AMxxBSOtl9LEYrYl4Ix0MyS2cf1MY+TuPRo81Sj+wTSLDzdkhRZf4jqVCyuKSR
iI1WoF6iszbIMj/k1WvMXf/s/6vbO+awpv8FDMgILCJIH7CB2xMJ+KVcjauTgME9
agS1FmtymZgEpa2cNpW4JiTEdL7zzF4bS/ugq4M5xhQr9+ymPLCrgZnwvsndjfY8
Uvy6UySL7OQ74j7l9MupHgf6CIdt3iHKanqwdZv+eHTbCTjWe2aG60nF1EvEqcRt
c/yn7A2rJGRTEDrHMYnY/AoPkqTt6jPb8YeKEiB6WnRcE1fS6Uo8TYo6Cb30niVU
3c/oHjMTuDMaPfErU8FC9nikzwbE0N2W8aMWfRYHOc2RTc7QDKfRNFWXq8xIcogq
TRkBU0Voa7NTIaugYbJSSey6iWhoSwDeQGUzRU/EZHIai2jngIG9jN52ovkvHqrA
1cAoMcvgcFWdAHABBPYRzfR3A53S7DKnExT+rLiM9FAi1c2FIOxxncH/aR8mpkLG
pmlTaFBt/gUjKYmeDDC/xCulXdzW8ElztmKBJwUHYRb52uywP2v4ARWrXPoSvvUD
rcED9TkEXcu4/XP+7LLWOS1qMO0HxILTlW7CphiM8D5F4swzOGG0mZ1rSmqGSn4N
jd3iIsjophqQP2AEN9ogUFOe979I5wNX0JJWABMjmzr7wGXKFQhrTX6Zm7EfsOdm
7k7fg0mGWuYg4gwvU+QXrO4LZFtVQRuVb9GYbvgiFWchNNe64FdL+daVLV4/GsKb
qW8lLZtn7oqy37U5ZJeXVQv0wpDaZKzKrrcY9UjbkoXHskmVKKe0ZxCqSlWSoFZz
nML/lj5agj143FIx3M89Se87EqR7/vzWbUgbI96HMycc8psU86ZycJIAwAv6Ban9
/GGH2JJRrSa9hbxTuPQWmsB+76QzuI3ZAJoQCP50W37htI3jqF2FSSmymvZ/0o0W
5m9RK0HIYWxoH+YSmNt6teQ8WcQFnBJS/yFqT3c8UF48Drrw/FeXNMVl6phpQtIe
THtYWZtW669YDQ7w9r4ZpNfN7MsFQJYjlXGgN3saN8DKyAwIZIwz95XUPyqfrJ7L
nLmJ4O2smQYIbiph04Oc4WcoGr+qXHVMvLtbqdAH5LCciXTCtfGg3UgBZp3MVn+k
db7/W4PUkyOSFZ24G6WrLRSWF3NPRzSB5algplT688gg2rqT7Acj889IN8aZrXpc
vwGk4rNCXekuPb3r3FUjpUfyi5gLbZ9V13acim75u++eKNnhlptUSNWAPTJegQX8
d2I3YAafPiCUcbLMepEczdc63OhzbUWehns5wEbVJg3FcsJ1IGwJ0nGUSFQvW6i0
y+n45HCjs0YdR1lHiK6dA7NEIHZ+P9UQpqQhhzkoCqn7nltwi8nLH19QIlPc/V4Y
ODQfAWiIOsPtruWjULWzvyrAPHK/rGOfEkgl64Uyzoo/AiinE9bOOA3ZrzoVPKy8
lt2REf6GD96qAy8YV9RfxHWIvJ7hYVyyjvinjwZ5F0+J4vmAAzLx9IaXL5P1Hk6y
efvvX6ICLjyT8rNuw/tLakVGR4tG+5xqj/H1gVT392jgMsugVMFPEOXYkqNILin/
UkTbNExxvceh0mE/PqQNZV+XIi4Eu0NdD/2qYErirrxXWmoaWY29WSOcQshlXoDC
mTHZ3wGjLAO8jJ3cAMVqkDZTrUp3hCStA3Md/P90/fzXSlmhMYSZt99/HBZRKKSw
4qHYCWmJoRPXvuxgtQu5pIQx3VgGxSF1s4T4mrxf6WQxgbg+TjXyNqcSg9JsuV71
oP7zMvSraiImI7uvIO8uO0lXvyja7DyvruCJCyG++KVaYFlQ7u5NYKa8jWBFbKt0
bwl44dHVWYeB3iNZqDWwEXOJVWr8fhdUTfgbis+esgUQInBBI7CoPO8Id/pf4sTs
Tahbl50OvnHZFwOh6vfNNfIUeQOYZkv9yIDKVWDmLsB3hp8eJfqIkwNZbfiXsiTD
n1KoicaWTA76SHGrppV9qdDSIILX0C2vQdWiP7h2OX2WiNXHqg2hJJkSEt5b7WU6
ZO/WQ1zsPEQSpccOizPmcUuFenuZiUBghN3eYgYe1lwNddfCVJyZF3SYyPMl1VMQ
gNlEc7YrRCBZwIWRZ3y6SH3SHueAz/UpxAdVrpuxfhj3cFAV9ypUq5W/GAzSCoNr
hK/rxaqirqN8mZ/Tf8EUfBBPoy7Rd0d4rVy/gscJjNJu23t+y4UcuvuBkXoFoMME
hKrIqLfZtD9zwxYpOuQfhO+ie4qqoooIpOIO00mGOwl559YBPksKB8Y6n/h92rvO
7bQaa9hu8XRDWjRh0wiYwSWlUqBF+DTwiLc6owepC/bb3gc3iSXrHcbBY2mAEMAU
XWA1X7mOkSDMf+QVXM3U/UxW8oGcQ7iNfaNpTfv4w3/5v1yLmPGHqchk96walnd5
izpwQhqcaVNo9cHoaE+e1mFQvbNubxnJN13wQi41Xy0Ct8+tmC1YG8bPSvia0RnT
2tLiIo1eVf9bfp+W6fNJBZHzKErpSnYOuWlgPusIDWLCciez5JzkgpMlKTwif6Zr
jsXP6zvXoOcjnuvNMZVx5sXDlaMDAJBtwFqIOhy30rQqV6tH9aeYPPVlzQVRHb4P
GBhKuQCr19vxSDKKltVJdaGWHd4ytdSRHqS82o9FW2cXZhQE5djkIXt28P71t1Tw
a9bXF2E558BPOQXFUJ8onIdnKt1M6Hf6iDNelUZA6qyftl6n8ipNp2MsVakf510k
zVgdtKVR8IFaIJCunlNg3YaBd3QrOaZk4ymMyvIj0EWPYq9HvGWtmFrJeuWdDm6d
JfeZe17rCGu0OkkurJ1EW1jdHsmUQnl3EMgvOL31a8vq4OfPIjQW50EIjRx1oMdR
2FsLVWgtcAto9yYtY/JjF0GlEwXSok8y44BdOX91ut68iKkvdkKyU/WJuUcHd5nz
UVJW+D6pGrZG8vtueVXDoedJdwYXX2qzTRLN/xl1AgCQ/DPdLBh4ac79g+W37QCc
4kA1p195FAEbj+EO1Fb8k4ne3A2W5PgnrH0X8x0MMcPheXm/iBFC+zqeiJune7mD
GZaEgxwtkg43b5Gn6laBQIpinIMBfr3LEjbhQ+1FK3UdYJEdLE9GPlQpOIVy2nfl
E2tEEZlmnhcwqvdR+T7bSjEpv8gDK0Xdbg5ok1e+Zd+fWXkhavCtuWm3P1OzjhLR
SJGeMlCjxRudqAWjSqEFaQfkolfOTWKHbQy0oo13RGT9Y/NKsF1OG0Fb+PxDtr4I
cUGtrw52WFDr/x8ryKGqGeRr+uIFd2qrxPd7VJPVKIF9x3iZXsF5PU/36pYSnt15
MiKCqTr8q0lh7VqVNRyatFHF2C9qZmvVByX8WDCP1ggl8XP+TXUxX6WX+hyyxhg1
YkPqJegR0VgsIFuJxhWUPAsw7RFCUnN9uIkJlwB0UWmx+wKWJ8FzYyDNhVvY3xif
PmQZ7RGCC/G1Nv2w9IsSc7Lyzddxj7GVBHAXn00NRw8i/MKpKasJ6/5r1j/6vVWY
PMlIja/Mg2BrSkd3Jz7sgF4bzQlBzGi1neX5P86Nsz5UAnPmETwI+oTxknwxyXU2
I/CO4Phgljx6ZJ1ivwsZSJ16+deqB3W1YtLgzOO24ih/575k4m5W8gtsHrjGmrOo
WDNsj+VDi7lxOGgkSMAQCX8awXUwaCqsS7sn/zxZPgUSI/bYEQ/xt7Xz1abBqsry
YYzfFNttJLAF71YpfqvfUQw3jL6zdCbkJPpZ+9bW6GhXXTnj8skvCFxQbpO8ces/
JqTIwab4hbnHDJFzAa0wLoomGlFz7R8OG22zsi5ZDMnXSL3HRi6Z13IiLTUEsXzm
P1YRB6a3JpsGkW3yhdHlaLQchv4dVvFaujgAmP7Xns51iqlRoX/VXcK1242wyjJo
NlPI95arHT2O3deRSHfFDK9kX35I+oCn06C296xLvgJqCDOB+ECc7CEbyqlfcv/y
pCYbcky3CMYrK0+zrzuJAcWpXPAFqwDHdOWj27gfKj2PSACOz+/8f3R/sVIMcHkv
A07Uyi7IiJ5BevoSNvTpr0cSqaUNVyjWTT3ZXKtLh7GW/HKKv7nR0mqFXgDEFGnh
7bE88AlUWSODvLE1StMldfpxHlr+3brdcr1rYnFhwq+TpWKx2yVf9D7WnmbfFjPw
Uh03Q5EGejMSYElt9eyqVhh7wLE6by44DAniWh0LcPipaYx6WfrYapwoCcjWIhLk
ECKAJlK2JkrqclyOxnFgncmsVywmn5FRxg01NnQKNiYBYk/6xngR8B3eGSbKNgSt
xYbxqDWYGajq0p9HXwkNK7OuSY0302EgY8iSGLfhtyayOE6Lc/WPhnEiPVHZGDTN
V7tfrZhj9+/ZOpivAb1MCdN4faGqjap9iQZNBjPX/bxhbjZtvZPhvC8+at14c71E
HNeubIYGyzVT1ZiZyZ2S+oodFq1gaTETjZpVByYvVgO0Lc9zKPW8B9TaZf9RQGgu
4U8FJf4LIqL/bMKf5JnCH7BBee1ZYw5+8QD78oqnNYVzy55YizvZmKisTo6hL1Gc
qFbi3tZIlkntrojCDwZIM9rlRm67VDbsaI0HniacJSCyaqzEYg4vjh2IDUZop0kV
PvriZGaFJ1FJObXmlQTGLi+npKlMIgrAk74kXw2RscpwOxLyx9+h5JWnT4rBSPg5
OgYfPiQ2uHulZrt/JyKmsWlIJwEIqFJqSicZKrsqPczbe/mFwGD8P3/k9DhBDP6n
vo1UM3pNCiBeYbYP+bkvJzFXhMsQtdirojCYjwhgGYxnOsfM5muGvjpu6c8AMjCk
26/EADZhs3DgwDmfDufS9QdYfz0q86s77iL9zowgrA2Wx47UI0EVJLFcIle6RXBh
ZOocPbUzMV5bN/PmAnAH6avpLYwn5QpaNYvbeZliB7O7k8FoYnN5swRAmjM9iuuF
inHonJ0c/p1gdtoEAKGP9BZTZRTTMKC/EpzjS9UyBHKzXB5wyfvNlYtsQMkY38sR
DNAG2Cn+LHn8u/Rxhf1VEE+JHeEbN6TX6ROu3Ei3r4hreg6fRyZfwKhqM2YwfB38
PTxNpe8GQmjX6B3VbdvlF3GOzJFJ/fVsrPgV+Mk2TvCg0YmA9Gka7E9XklaOJOBg
BM28bFRdGKD+eey0MxM8d5TEg628Q9lJ9Hn04vxIlHZ/MUp6Cv66umF0Ca/z92St
E6AY3JbeAMm88wFKIvj//6qEvx2bYeeA3bM3LLqiEo/CbqlLq47H7Wy0KkxmyMNz
ssf9xRBOW2XfAyZ2zsaHmzX2q4Tw+O7c0Kfi8qsCSnatRZFU/7eXDR6/j06Tg2LW
sLYDujy7sTMJvrLEhTdLBTLj3DyIDKDxWOVJaC2bCuwbtFu3q5TyijcNEjK9YbAv
OxuqRaDlCXMkPy2UjmGu/SghZdXAzhB1IAxUX4aSapZHBpwJj0B4hRTHR4CPM4Xd
SUkc0tPNu0M0Qh5FLkRxuoHV+1Wc4tnky0IpNboKr7zYX+XA6tfUcfRExE4gTJS2
XN0Bg/DaMsUJPXpStl451mfeCIkH/TwxYIei60Ci8E2inYUCS1+hU5aLlbqyk1I3
H2OPklHavNScsQVV4pL3IoIM0qcbQho35Fo2h8vROxUDWXLStbobY1JLIXBTqtCK
JUDexdnoy1dmQnflAyO6l1CVc2ttAmn28Acp9JrUkLpueK4/cLmTBKbZRxlcfPQa
i8NVuwSS2CodGvVoeu08phI/p39F6NubGJX6Awh7GvUThkVtjGUrNIElJu8OHjd3
pA0miH4uF85S4vPbjSswO9nERmjLJ//c2VG/Z7D+QKTE4Jd5yjtpf36cRErOhUMD
AhjDP7WaO8NvikQcGQSuGZtCFy9wmkr2wwxn4JsDaPhXdl+eV+cctFxq2j+SL29q
XP/3lIl0NIZwY3llsncVAKvh5jksZ4lU5DGRpKRng/kKs+OaaBAR1m0rqTpSiBIU
phoxe1JxHLmwHPCPw+zvT0AUebL4mU417sL3mXmWyOw/C444KOsgdmrBLFe7f91k
yHRIfrGZiwFXZxZMe1nJKChSg16LdBulW3By1wXe429bXZt3qlphYj9Y0BUG0Lmr
oIxfxovc75B8dUDgIxzYKy4+fqaVHWSuFXYWEtEKaYNDzPcXp2c51xTc9v6sf5Uc
yVoLi2LeXXxboRN16KiimMlN/LazZXp/01XJ1/mclZohcIE9IdpJNAoTBTEDIS1H
XU9dLDwdnyx5skMQ3ps+I5BcPGfV0D+FzDG874ofKy+U69v2VWw/pA3+CA5RmVhU
pJY+FuLb6vn+n60fDjJ3EQ5mpWK8kR6bNFqXuj5+4ecR7pxZXuJ2NxjuuCHo/XxO
JDn2WL1R6ayCi7DCIy1gxRh08rSkmtVDl7s9rMCJoiWt95AsVVhCaxmJRJJDeO8E
7jYRh641h2FuIuN2sHKivkE5orrM4syuPl3KL0xWB+KDGhZhfiVESV9NAjm7edKx
wOELs4osxVG8me5cv0zkEr/OZ1iXHyhZajWn4HTzNJ53+MI4G9f1obeolFqIb6c9
I6l8lOAf28ZCQxkWka3RZSPn95ugVhn1NcgebAzlNMA3pCXLU0zOzNyVZLjQMnvV
WHylU8Yh+ocKNh+LkGEntT644rlnR3N8uE/1IL7oa9BB6EtqD8PpCkseft6eJ7ko
NSkhRriyNNquZ1Bgy42YqMl6oX2MOy33vfXv1YfBmD14dzZUmkqGntmAnSPbfhzP
Rr/YfYGsKgFPfaY/zqlqyAiBGKDqkAlykyihrrpVV5Cd1ZmJNsezHZKwda93hJtA
6q4JUuuDz7kVUf1uLx9sowuHu447M2iE78GcsB6lHVvEQk1CcisqVA34+SJkyooM
TKtZ2Sg16PIKQiePHF/aOi6/60M48dtj1n63GjdZYe+VwBStJlwpUriTB01B5Qs2
C1xh8VVvS/lvkEgP1MELI/VcM+1/h1k1BfTcFzcYaMG2PE3e1QiLhgn/CRlyzNXx
GVFR5sGC2/mtAHHXwxGKspAK00hW88z3AEoBhwG1o7N4/NM5pC3n4CuEjofKD5OP
cOzEdDPfn5Ov6mb5i9J4+qlgBXs3HAYD8/0IWQrZIPCFOX74cTBxGckgzypSQx8W
zkKwTOhw7PxUc5bIxg9nR64+FW/gIXsdgai3jFxA8zzl2OETH3gyR1CZmOPDiFaH
fzROd6AxRGaPdPW93H6JKnF/5offiLmKBQQtzrueF/V3SjF46VhYwFsGDCqvh/9L
EzN4/aaBGN8K7et2mSY8FRGmKpHpb25tIvSRb1NKIVkq6AgUXYvvI5Mws6/YJTqm
TgV82elFMzPJWwTN6NwVlbydKbe7MorCPwTGsutd8Ymolo+DgonPYRPdb/BfSRPJ
3KX6sDdyjPrwB7N9grVgR8xO+yRzHsse63IZBnEGo0Qw6jf3+UFNFOQhP3VEkNSj
EwSNnNCYAR7vUqpkeLwBZ5lqIJ9GKKLyQ2B16EVZv1bEewcW2XBXXPIR1piA4wpe
XqcoFjxyg9mCXImsln/ku2T1/oNAH2h4es7ENdI0ZuQkLU9uRoojLdWQ8f7yP0gg
ZWC1XneXSrSnAdOJ9qHN8JOilvMbHWzGVUA3tPvDtHB21l4Yj+dW5sR8ccM0coN9
ufLcHcm200+bahHQgwFT6UaxZM2CxOcRABYOc74xQ7Nxlr7fqvo6PoXLTMLHf1yi
K/xJhscDQ9PI7u7TN7TyaLkGOOTtjnxAMapgDAkmmZeIrSxLy62/YaHm5Aki7jnb
jy84PRM6nk16ZxOoMHuTsUdgAt5YpAj5mpV7uPGKcR/yc3ZK+X0mm+uZ6QSBel7S
EUpp/yLwhFcG+0n+efJy6lsfqt1vuhvKlDSjCXyqYK0fq0z6F/B1AHvD4rqfmCGC
QzlvN4G+P9PD2PD1XuURBbkks0ajy6veeK8kHEYY5TiFrx+CIRHLApBOuKE1hARC
Q5MTqjgNpFmdsj3ZuPuHXCv6QElJL10dFyAriVm4p3sYzBbLCdA25AXynxhnjHkP
ytTxBeggzwKELZaJw4yveF2DMvz+P+JZS80P1x6GTtsoHXGi7Z7WBcXcz8nk7IsG
Az0F5OU8+SmWmfDn7LIZyTQ5DMbrxTcuajVusdh7377cIFYthMwnF3FMc8vdVazg
jlUqXqdxnQJCX2IU7BoQH8bJW+XNip1tsO5/Dnv0MwXRMTy2CiJREJ86lN9bWxz2
LBBTOqPIAG3LsmiMWwXEkal4eR4voc8j8b5HYYU6XfFE+utxMpLt7GFoIbIjNz8q
AA9OQQSvMi0Yd6OtCF4OIrGHUiU2H7qjJEYDXjYuk5y31aKrIJhwCa6oHYTYelyN
GO3RWpkJOdBuQ1jHhYI5Ensyu47GUi1iK/loLdvZODRHwuCDShKZ56iiboZvYNd3
kT0ksOjZN0QOf3ly7JzZ/NHTvnyf0xifWR/v0tJ2Y248GJyFfdMysVQRnf5zUDE6
g3+Iud8CswpB7G59nN6PZoa86OHu6tMeZkiEsnxdsIkCqG4JiVxRx1/IK7fmrEvB
BCnLQTsMrXVU7uu0nXOLy98PfldIHcBGjHcJxg8QYOTlL0n+8y9mGYdWiXSTvv+m
qQMv/u+1eLUZ68GVioj9+gTwyyIF+JmfRo1va+qNCNQwGA/dPrcjZNun54EbGW7W
o8XxxuHqKrl04mSsgh9ObuOc72j5pSv8u0B9G7lCmymBMiiJlF9qGWvtbLJvHGfl
Uzg6gPwITgXKqHyU2P7MvSHHHypA7xbkkQ3Zo2YW7nmVpz9jQ3RMmo35vR8k/+8L
wDNztoeEvAQg8YpTz7wD8XNxtqWD83HKXahoQgom+luIZqtX9sZtJHlZP1jxYrD3
N1XMy5PlmHPUS5b7nJO5V5JgzWkRG/YvcVZO4R/qI7l0PBBgg4XBh4VwTH6R/XsT
sCW4rGv85Tn1zxLOIem/2PD7j4BMnR2aohE8I2aFH2DxcmwI73GnlZ6fvBicKump
7Z5IvsLr9Sn3U0LADl8Mhr9K7CaGTsZ30YDAhG35/L+XyBMemX/ppR7d9XEWBr9V
+gor8fZqTWGmG5oo380P9UVfrkWRQW/66kGET9NgPQRl/1G+dZMCk8dhYz957ADP
JzneUxBAA6lkWbIZfyfl0b92L+8LHqrVRFGVRxEcq5nOP2m6Fxxhl19b83rF/U/3
YkxJpu5L7iJ+COGHDPARm5rAE7IURvzJEjR3Xi4QI0okG3ab0v+y6+bRsHhNUxw/
Kvd7XUjGh9ReH+yfBFna9LGJg/L1d8QvdnnlHSbP6HFPnQRHs9TZRpYquY2Ic2j2
0/p2c+qvJFkIUk2jWWehGTA/l+l6VNn8L3M0MXUErqfcRn9CYbJDLj/qkD19SpTw
H+Q10APoHNGwgdE/IaCI6wE+WB5mgTEI3z4EC1R4AlLni5/LEg148wYTQugfi+34
wEQucCBGj5ahZYGUPeGoqy1lXINhmefSb/Brfsy6skHcGpYrKHYNuNfedGobZ5hh
8i/7csJ0tuZm+5mQT5NG6kTkb8Jkj9C/hbdiN4djYiubzEeRxDpY0rLBf3y7RPYb
EMIqpp85gNKczxJX9L7IbMizD6povWs4qSx7j9iYxSuSDAQUGOWM8GNvuSJwPJhs
vlhjTW3NoH+i7IkmrmfUeTo16vzLKY6pKu3q0nUFXi25cuH0SLQeXhOR0/o59fv2
a4jcAJGgUJbbvBnEJp0QzSsYSIENmgFtT8fhBxr6f2/aMrIm+8GuWxbrI7JjqYbl
nVnSA9BBexG6nmb+KtfKA+thio01ILbNh72LMXwCWL+Ozf+wcMS6jYt4PeMVcsYV
ij3KwaPkyB4jKctrebhFM/yvd0qECz7V1lgq0FDBf/sHxAxvQVd+cliJ2LGM4t0+
QyNT7XOYf1fAMHvxrDifDr750QOylfgfNvkz99+HOug94yCif3qdRS26TaU5yFsC
/uqcioNHMd4CK0xl7x+P8Y6rhzHxtw82EL5EZzaE1e78Z+EDx5q400/8rl1Xrgfs
UmUZMD4qxEZPbW0nXCN0Yma5XGNojnw2Eb/lAPQzBbCOZ1KpGPgDoNr47rEWLlps
bFtHsvm7rOycOOP98SrP2JSlc4Te9PEj3x4R8/Rcf9BKcDG1a5RBLVgtGjDhH6bP
C0w+xOcf2c5lKU87yQAZR0MApYcjQEcl9yzfR+Bf0xcYOfWwww/ACKDGqXebabyg
Ytqlvc/juunrhFZk+hW1sLazmeitoS5QgCYGMBYBZ4x720F+e2OgM89GKcz1YNKC
eVRnSMG4gIIhVxiGdfEk+XCAy8zpr4ht4mQA8efHHZ5wVPyLM4Pw0tf717M8mjgz
0Ony6x/XtI2KcWVOIqL4ifRgOa4fas+SuqlkjOBG9SClBzp6SlZsj9OdAQac6h/Y
mHEFzUo1Zyv4FIp3kHp9QE0u4Zg1Ij8rcDWqm1JN4BQILPfVhIf2JKBwmLULQw5I
/bA9Nrm5dJ6ipkW3xRODC6dkjZhz41nnLnC8r+jqwQl9+4ESfiCpbh65HltyO7cR
/YANoo0k6Vj71DLza0KsLb9pfny+06q/ct7I5zEkH7vKph8e7zR5Yvol4Qrb38Fn
0+BPawSR+5/0eDre5X28FJBsDroK+MrroCdleDFAI+bAOb/GdGe0Y5xsS0lTecI/
qFU8rKpqbBx+K9XBGDtpA8WvVORJQf2BR5FWTyh7mi1GgMyywXITvGr+uQ/MC/nG
/mJ6unPxIgK8LbEIo23EeMTCOmP+28UOVvKRL7JGFrviiJxeGenKM16nomJ58vfY
1OJlvPDIqwSCtFZWe3MsBhW61oM+klxm9H8lMmVDHfJHbFboRoCijuyPlczEksTv
gGsBsvshAC9z4PZskhygFbkIuVPyMq9BfBUfW/diWnPexZptRzA0WJ2YUNXOCL6f
1BeF4n/eO+lY47K/5qc3gt7nCGhgzgq6G6Zr0Iu8F1JHLLbdYGawNl9peL6Hm3cM
psv0LF/0ebzZCTsq5yrLCMeKx/eACF6n/DRFtJwUf9VzdSyj96GdaUvWSbQuo+qS
PtGn/CgxeVeUGokvoHo/9JLRYNXedQ2wEeAC++1d8omSCnauSNrVAFOiaWiTh3Jx
WdcaVQLxGBnjmUxLDIYJ6M0IE58IpnOqdnUNNg/mdUyTTc2Z7u73nzQ5OZAU7oKc
sfQh8v5/QI/ZGd9N4vvSRovEGGXbRj1lZ1hwvzjEm6aDnKodnXfkV+mJzzuFYQFr
iN/59uQI53rkdcbPPgeKTjsMlzY66sULJeHVu+WiaAn3YrMs9DdMViUDxk4ka61J
Vd+UDNvNL3NNASrJAsF+LuAt91810c+creYGipB0gqMRBpPZUcUlTOqCvBz6Fc7n
J8stAPHh21PKLG9ONrVIdYom2tX/E/jRQwoQGvpukeKsHhmgqIzJ4TMproNEBaqC
wMzb2xJAfuHIHjLLRhqzr+jfgicpZvhqdGcTshANZJwOYsezMHjHMF8dJBjlXb3R
A77LI9uXfREDbJzq1jWhkvn4wO2iUpMegDsNd1/ZgDHbr07Y8svuv+wVsQ7OVd8h
Ue/6S6qb7YboNgjElGXE8CmOjjnuBUMQpFObOzNCxDM2puU9RYUsXApPfq7nPgZO
j1yplV4hPQlKIRTgQQguJ9EWmtCO30oeeKb3mRhiyr6Nukp0MuPfd7kat+z8Mo6n
HNmqfd1MxA5rtF5GrK+Eah/0GbLaOAGgGiPOebtnozW8Y5UDvewfpEdhLwP2LomR
HjaxcDOwMtnR9Rdgn3JxJLb9xE3YWfxQTHx2ho5MkeiT+MKgxeZYpGmEgQLMGZaq
dtZ+4M1PfgJLl7GRpsKXs1SWjDanFf8QKRiFHuLGvsNZc9B0889Nadpdrnvpi09s
6s2HvuhPAqeXQTRHOgswhSy0HCZc4nHrAZl0frgy/U6uyjSad9js4K9bdiAGa7iD
sG4QVSV5nqhTSTEqy6avXwDe8gVwreXWO33FAvsTF76apmupXGvq0rghJaz2XOCE
uXkPz6BDimhdZ5AVzu5QEHBel8U3XswyMrUqfLfJ2yotzPJIDLRGkX5QDbSWa8NJ
ZadXVrHh1AHY6DmNXmd7d+8TICEUrR97Go2WWCnqDrWqOl7w/0JeoYzrm/r+Zqbz
CxezpPcMLV2q0QdGxIxEWYJhd/g/zrMxCbQlbhqwuZAe0u1rkqsMCUxoYtN2p9cL
hK7fz1yZK10N1bGrUWk5oqi6VE4+7vIadXFVAfgxV24JvhMAe+58kkhKCD1lw6CS
++CorSALtHXjxRlM6OaiDv1K6muTyKw2YQMbnJnceqfs/ZDOyrQgeqUFr71jwXYi
0w9pR/5DcqkYs3vgB8yZGi43Nn9QDTb6RLJKVlzsrssc7pCnpTKyD3ioNDu0qRsR
/GgBt9fGs+AbF0Jp7GWkdJy0r9z0JOyMFhmKy/mUjL3ubW0hlIOPhbenRhsfC2jZ
0rtMHH8K0wplS9OA5h8RELf0VNFKFIPMHsx74InpkwRGRMUuAEwRDAUC0HcsK+60
X94RvdriIHP5JJFjt4jXnqNhc/wR2kxghGWmUErdqVhCsCFcm4wyGB3emONKmudY
EOZxDz/smC6wtmjBxseitoKRdvqAUC+lEFJ8ZiGwQv5invUu9xalobfdw8XWO1BN
EBC4rwh/oACb7Jn5ZEBESSPOR4TFpSI2wYI2E2UUKmAiW6vDPsmVwxePqg24vlhj
Ue2ZGY0GJVZn8FynDb+qqwEdOI5Dhaf7Q0we7WV72cOMhtHhB8IInujw7s/ImtJE
Tgz6eNC04MO9S1JiHpH7lwN9Qqq8nFkb+6f97MK7uRWDjR/gLqPy4PX6kPl+eX3I
KGVF4YwsYoJskF/S3Itry3KM9xDXs3ELOcJ3MTyu8cgRj4UK2BVzM5f2Rri1teGG
RvKSrJFL1FTwMDWl+5Z5xAnLjJpL6G72714V40dp/qCdV8ughNCakLUZUGcru9HM
VMaz09+OzN8YkVDVVUojXAbTIHYq45YrW/YQLMBY1n9JyEgzcIGYNjG/qffOLxjV
81iqbM2b32vCMsrYpjgJiie66c2nDFvt9Z+Z6ueg5d8tk7lky8eEcENJnTcKpBkz
rzaiLwD++Nw0oMDtFSQh2u2oj8z20vfIC6MBoNqbO3lns0XnjJAwKdjnPCLZCwDk
v4gCZuJ8imc6WSt5ptO6xVNV+UYKZQ08d5ACSk/3xryOyO+0pprybWT3esvbeK06
riqQreUhUbcavVNKL5XGlDGEXG5L++OHKCeDR815mRNek2Jr1oXz/DTQszL1ojWG
LzABwE/goiawWJtNEkt6DPeoGjG3hRBOKutRsdQtKWjhM+H8sjIr9sV+ZI2GFoJy
3I8FfvmcBSSuzQOp+KzJBgSbHzkG0rnRnxMQO9sIZ6/oqDiB34W0OEzuf/NUTPFX
MrYWlWSXezdsfj7a2SkPrvvxZulX/TfKmMw5cQdBSbis6aWN2zV2acmBUfjZqy5M
+6E1EqRLZBDRvI4Sd8MXnGvCpYgyFh4O3is4DuL+kXhEM7q2UYxYOAFaEslG38Po
YBmmvMyycWqHjZfxwakdU/iYV+YziSMJxWqk2HKNAt3pakbB5jU3+NHVKRCdRyQJ
2+yYxLbtxW8oNyM7yPjy8iY+wWSxhHV4oq4L5WN/14eJke4RMzbl1xuoV9Szj/tH
yKaAJuUIpj77CwWWfKvhMeeT9wEzHZXQf0++vztUbiwDeuBEMNZbrC4XcvzcoHWj
ab292ny8wWob0xb1v0+kW5yRre3WdLSbE7+2R+yk6tO089NabCWRHwi7sGfDusFs
alhRsFiqZAXamuBZIL31MfpHbzc3cUvadzgGr/66SOMgQBPJ6dabo5WVHcH//rmp
90t/EIxVWHb0kY+c9y+QdNDP5tjR13MeWeHheLvl4k1TLrxGiZ6TpWUh3e46ThZh
oP5vP3hm0tyzWdiLxbTSzt1XrAuBLetaRPTKOjS7Gy3OYFQlwsiZ4kq0uxPREkFu
CbAsR9vm+Lp9Fcrvq+4nlyXAWJyBjmLE8EZNQOoWUY3tq1h+uP4BW+b7J/ZD/pu7
aPDXaA4QKu8BA9qgUkMOxi3CBIPXAd+tpDJ26FIDgI6Er6rWRNFKVylYG84nVbO3
x9YQgHFlcK6TFiRYyVQrx5VEPMqy6qMiG+qD8yRYnL4yEhICCHlrNHww1xNoaivI
6xW0u5r98teawpReyyer+LOQ34aOoUs0ro4AeB2DbC8Kj+ZyE1l7ys+vj7xt0j1O
YoAeoWBxGHeMstYfFZVP/LFT8UjKffEiQTwqsgwZ/97hOn8gl1RBd0/Zn6FZ70Mq
QdpK6cVW1ZyK4v+ptdXx1VftlBdRXkH3MSD9a99oKaWSLUBHmeLNE8iAtxcKIiij
x2V0/cMIxeWdWZk/qdVyIU7ii5tVKgXqmGaPAoAmVF/TlNXF4lGJdKara20Oem8r
c4H95z35n5g/VuLYBprVEuzsknh2YkYDP1aLhS8F1XA1jnLGnzMFWnUzVO05HqOX
4LqHYeg4B7zB+IU4i9qMWtK2ULHubfciY/L8rJgRoz0uPDmYA9hMwxwtcehg/Eb8
wIPQRSxyOjAxiytvVXk7Eo7x8PS4z2IIVHYx94MNqJCciafCg71d48abc0nTF5wG
AM3WlpHwcqWww9BV2Vc9g8mQ9VArr8DvveMVHr5gU5R01ufstez8X/9lpZDo41uS
PcinxJeRsiKN8Q271HN9ouX9YAGD9yERWf2yP+Oq54jbxbGYn+wEDDD4SVL6zaAZ
uvY4xDd1tkvFakse6gyUoI90Hht15p80/yrr+o6gAvhgOr8TInayPJQ0rMem7qEM
STHk4wQjf9bRAVU9iw68axqXU7prPXD2eoAR7j85SAdjzhArhaGaSsFn+GNK72y6
okMDai93GO/1nNm/+kXtYLzlRACaKrnb/h2W8JjPbfKt6IX4i76m0tTCbO6hwF5V
YDVU4uSD+vHrQVUyiFi2LA9g39uSCOS7KrK2Ws6gLqpiWj5vl9btuQE9h9haUqLP
AAIb12immiSGLxEBaXnPSyqj0cLLNVO9ZQcry2G4uf2rqWxgCFjZsZuWM/hBbnzL
CjFRxz9f8amRZr3BSikGwC6OdN0bDZ/1PipJ7asbv0htR0rQmpKu1GAW5GIOWsot
8Nqimr2TUcja7hpxAyoM+arzc3h4BzMr2MPigFtOuazZcPZ+tI6eWyMv8FG37wHu
2XE7VjaPzfSW7nw6LApikOnSQ/qUIVfFYwafubClqpJa7tf6h/9qw5AMQuJBsUER
rcdt7+0Dqx16dKfavM215usyFged0nl5TpE/2AIJ77sRQV1Ljo5pJdJFGpbu1mO/
ZvIifVbZTJiB0asO2h2dNyu4/9q96W5Hp7cq+vu4HqshyV7DTZQ2DgFh3TEVxUCY
9VmrT9C/Kw3QUR7HwN5V4eBLIrB4fJfxjn3WnXT2N+/jdSCq0v+OJHC2RxlfkF3j
/hpcLxA6xrJPCyA7CzRMe6RGNDAC2GEiAeBs2ffGHfGkUIonnqBMtedP2M5UayRB
C0fvSu085gfoGKgisA8XUyK/VbpM0YV53ZIywcGty1xzbgUV9wKJej668Vf91AOQ
e9FGCmviVC9AEyWLMd7iqqS44FRgeZU0GSU77Q4IT5qnzk0NGyhMXYi7byQ7iNZD
L4dPn2J3XFpgV6cw/ywRvW82lv+uLRC8VVPlAvhKHkibiUsuk9FFojA+wgb9wAgC
jbogsFVLMqA9JhlbGs66iHZvW/5JwB+FELszY+h+g7g=
`protect end_protected
