`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
SzsDvnDEvjFBbeEyt5VBOvEPx6xzX/yuBqF1KstSDrauDxArR4bq66IOU3l8EU2H
KUH0UoZhtRw9EkWpLTKgwPzzOxn+EupaHnnAA20r5mlnlGLAyz0xWcrMXAouBLQo
/gRJSUlJCtjpSJqGL02ni2SQ1qjgNIq2WR32DvN3S3cR+PEbeN2JsGdFBRRO1dO9
7ukiEBF5xpLRh5lhuLQDgLqsh89EtvTswNZbxaBBu2yqqRQLmBise+Qvx/PJapC2
HuFurnt5ch7iXYxmB7lunKACgXCHBfZLsbsNPjKd+/7ZehRtRguFySp/feSecfel
AWmwyyDwPZR7vCFtDGfl5A==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3008 )
`protect data_block
Kj5OKX89XdndOWP9Q22lqP8H80SHFHWVs75ZDaF0uv2zwLQFSOqOfFuWaXMoCv/A
9sXEf1xWC5xINkLVYzp7j8ct3EgrL4D1nf2Mn2Oxqf1UvOPIDRk3cZInAjyv4Skb
MRmq5Sl6LuUwlZQUK1uwa/KenaTUQdmtq5n6yvCWquhHviKU4rG9jfU4bLqHYkTn
9tMtU6H+3s5WiPDcyny/+UC/Wh05zahReBNcDee3XoCtE4JkBX1CVGjxUMWmyrqh
YLiWq6A8X2s/mtEEN/xBCs+8ESab6lrJvk1wKLyLlvllduBiu1CY1CUgALvF7Y5d
pc/F4qDk3eymUwMHGceRR939vsANzj39dOMeUn6BMy4VZ5cLXW6hEAwgS+6NeXgX
77T6cnb1/QqQZGBrJkECNUmjtArqBYATu4JMEiIiPzEylLLrRr/KV825kTeQk6vc
wSYaSo41l93uFwKAqylL8vu0l2eBl20z6lhY4+roF01maKSA6YjmG0OdiySHSsj4
xQ8Csd5EX27RjLUX+A2mhv6RmQB9kALspU0W+MxReBMyWj3yLtv7GnZzDJHrogl0
9qoq1ecVcY2zfajT+U8tmjICaaPMI3cekDHY5l2r41OZDOq8sYKRhLOT6pkSjy4Q
Bj7VLUoI6p2jehi8D3dCTjBQpyavjGfZGlbLeR5B8m7YOSoxKwUTZrdpIYKDhtXK
NB6vCTSwuOsYaVuW5878lJDc8zXDV3Xmi3oTmirn7trJjuf76wNUMyoHO2IxhM31
3fZoLs9j08C+xHwA+/U1beNPHa8xiISD/B4nkOuk5UC5rmFiVOYkBhmM9SXZ2hSd
j5g1CwELwx/ztjBo5oVKWReb0hPdGycVWeuuxaQYkyd8CplxGPIcbX/Fs/jGpcJC
oBZ8df8PTvxOxYuyKdyAGQZ/d+k89psLu7i6v8u5SFHDnyO7QHvNSwQiDiq6flp+
YbNRo336SvjF3F9kIgj2Q868oJrCciCGaUiKvzVbG3gTzWrLtioe+uRWyI9F7zJM
lTNzUIpbmc9nrNf5/a/0c0v9AwV3pay1z5wT/Z4SHmvhKTKydDGFftFZRbgFDTnq
dYtB4vczv4x++W/AmFY0dk5YEVdH2vGO1cq6/E0BtTXaiV6jCjO4kJp7v5h6NRDV
/V5LjjHQRaAa3GmjQpRwjfXLbvEui0oPUbWy5KMMAHmvF7XSPjGo8NoWlKBVslzT
fZSnGRCcbFP0AwO30fH3VuwuagQfFqIF9gVkldV5wkMVQn0XBXh2dTHxNK+8wq+7
NmlVhQw5Xzn/luYO3zvCJTUy1Df/0Lgxqohcw0beaqdxFBpKN/+W/uwQVdkJMWA2
TNDUK4IAhMePGduQLkrYO7QLDpjM2h4Pi7uhAfsrKXAdh0tZTJAkA+Rn7zn5dTAc
qdOVeaP7F4h1dcoVqciFDfNIiCbgT1fbcfQzDxsBbHb+te76PdG2yHXZ/VHEtbVh
xPRXMcnR3JaJHIbZqk3TXnw9nRkmC6RG2NxWSNKu2kFzewwKujw9y1rkTSl04DhN
rXcjDXkKHNWWShtljx5JOlrz8xlqIRLOCiwPHUwK7DJT26/BLBAZjw5OyQKWSFPk
TUA1ce9cKkMZvBBrIKrZ7/U83gi4ds0CCKWYR1FpSGs4qwDR7HNhxrKQS3Ymvg1J
8KZBJpZazdDSrY7UkOyn7T2msakTLnghP9ryGK6rC2hgCGkkdP1oQeobElKFB8VQ
o5aXrKVl6o7P9kNPluAObRekq8/gja9400aAH33+R9/0anZCBTdaZmNeqsBig3Eh
ZvOyH/82rXoCru/jHEveSw31sCsA73nIXaVSg1xXGrZI3aXlkw6v9foOiHoonttD
5jSvSc+Yq1dKZYjfWpqcKdNTrJstI/BEVlGpFalByc2uqLGZ4d8EFSpcGQ7+DCmf
qFB8+jdrJxDhIJ4pSI4/DUZjfFdhSR0Wh88kjmW49h2O2x2Ghsbo7brtFnfZcpNJ
0toSZAzMHT/ikJp1vqgvlCBQvezN5YRXcxf8gQeMuJ54xjemt2rpNa+fkIFVlsWc
fjt+3JuWQCLYPJlumLkr2CxdPrt5Fg1Pml8JTYhJVRVnFRoRDHIfzSNvthErfCai
wMRlma9flv4sYK3Cdv23MagklybZoexAzOoiAclBk264+Z3JSHrohbWcviNJqHKP
9ZjuBPBGYBAZFooJF91J74l2ost65u72MT7yDgQ/ij2XjZH7i4Dz/lPPncHM0Ntd
C6o3xKChp9SwIZLNjQEIhx22KEyN77HChabzutc9OYxUR06fdXPUzqFuG4RGn4hB
2d/r6psDPfC/hJgaXXOQiZoEHhKa1O8nZPWbuGLvf/uQ9Hnr6cD75nIOGQ/o6mcm
WHf3W0fx7A1OOC9xYp8FqNC8XUvQB+TY4OwnZbqs7VkJp6c9CEYlDsn2u8NVgRH0
XXYYfVNlZHVJkgNvDPAzaSOm6gS1x224Xpquya9tVqA3T1CfqT077WjVztqmW5QQ
JdQrf7zvxIhi4cH29sI10iuRy6BMZsQVefy0nVba9XERCdylxwlrVqDojfMXuEYW
PfYrOPABDENKsVpla2fy35iLy62T/S41k9fMcFig25lLwpiZamV5wi7cQzsyjwvn
eAqbYeifBr8YocdJWprOwl6gdFxLoVcqr4m3oTX9pYNFEBKB/iM1qDNac+g93WK0
K9pQKxiR/nEdNfX7nnIFj17tlEWz1IJlwd7kKutaYP83zc1vtveRt1uEeNdGfg+r
zRX/hjjPbFlMcq01TAHvIZFGMRR2QFe2wPIQygpYXNPk2kM1UxO+idBW1+6+ogpY
+kD/9lZ+ObcFqYbPocSahMDJKiX4tDk7f9DNhgQG0LdQxj8/VrnY39aKQZBb9JpZ
Tp8eysUXSKHELszUtL3R1NxG+X9NpgzGLTPz4lGu2oY11XKcgju7+Cu/C7877OqQ
+Y+9n2K81L1sguXxTxAMI8YY1vDICTXSwqB3bqzNdBEIDzhcRRu5lzgFFNJXJDup
qA6i+6FAoYVZ2kcXZMdDEDAbfhXP5WM1ISKFxEVt44kpJQISg9FSvBVk+BzZobY6
uOtWRvieSPo5ODPN0GiUn9h3E3VgzPkjk2uBXrbRJSfKyy2j0oRg6tq25k4XVoBV
i77X0YKUkyeamqAJraJll6zE/ugZc5ZVNJeUFf5ifqCpF3bBFR8tQtCoFU/EFw0n
YH/Kp2Z8Bj73yJkIcq+NhZJmbEIWnCY9/ukqkdq8XrqGqnM9cebwf2D+c/B1XL/V
rU7grtzZWImjhnAIg2Pyg4k13jg54GjhfrwVGcc580p+aGVfqNfBJMIl8E9lvM0C
xalM6wmoV5wwApAqEVZQLhqp0rISJb4jUnehHBjv0qsLBh/54eIpUtJxEqgV0703
pCeifot5VcAdzOqlzw0sKInsH+tpvb+ytBVYjaGTEO4DhZibydc7CXsrXieY7gyJ
yEojVw4YA0IB4FtVjSsCfUiM2TNhpC3DtiF2WaQTneTkH3XIIHuQ9zv8Lux2Mt3l
TEyoH8Nt5C5srgfad6fQQNUNcWbDFraJpURo3x7wfbap0x8ysl02x9SgAeYvh9Tb
JCmd0Jk4tsfbjfnnOS/CaToTdwlo6JnWfWhKrFRAHep9vhYp+vfcaPziaublNtnp
ZwUboVsLUhOesjbrCpCKF/ziOegUtTkBtCBnTyu7zT4fHrfuXONKlxeKIPNzsWH1
LeQabh0ic4QG4wDHhoDPkJbcdWbIkVOEj0tfE9LdEE/B5e/kPkeLU+Rkrqk4inVy
UcyY332rRy4K70GMCIJ9ZSBsNi8pvc1lNGJDPAD4nKF8/ZDULp5N5H2x+pP2hFf9
LmRDP9/V0SZHLre4js6DnK3DdeS5wQ+7osnLM+SwpTUR3uZV7w8Ap4d1pq1lxZdf
O6+8WOYGQa/QQr5HQNHC7slgQalaKZKgH4XXs5cPNWL+xh4edQgyVDHzPBPmLHho
GwCYkD/Er921CirDFfLV/aByVAn0NyJ8ZvjnROg9s4c=
`protect end_protected
