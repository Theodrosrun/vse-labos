`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
i6+tnaXxpWacdEB1e1Ix8RA0ulqylR8ldeZWi0ly5WsOmLDh/Qk+3RAfLy5zewq1
GqsevfFLDfgdMngtypvuCGSLhDc3kBKU0K80dTSWdtpUkeTkAtYFsPQMNu3K1eGM
TJQ1U5hVIbscEBNu8oUvmV6cAeK2bk2NTAQL7ZYEzik2wLCqjvgXt1vq/Ow76N82
IWEBMoXx0gAhYRWd0+i9qiJqpJj2LHG2PhwLvVyJvwT0ng7WISbWyrbfwXYfAEaG
VdvQfMp2l6jZtZ7yDxbY6bgbHkOwlfhxBbk3SfA+jHFsccLg1E0+gMUKe2RkbI/j
3q56MEMRRumzEe+u5VZcJg==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1952 )
`protect data_block
NV1MnMRh/4JDZ6tykdUO2a3lpaD9Ox3gwYU2AkQu1s/jrp1TJQED/C43Y4YB137S
XELvVP0ZFkV3yYzNd4S4SWLkd1dLZWZ6Zjqszhh0FeyTBs4e9FrmNEYo53xiwzRo
4tpNSUvSmVjZ4YKITxgDXbZC1P/sCfPPPafWmSv6t4Gv4KyQN2/zVm8EQDMu/zwj
seM/7G8w09hYLz79DzHTklOrakNY1IO66KrVNHtKTSrCm41IucZW/jUl4qTdWhwI
7pTE1y7bmYT6u1xIUxOBLCkgnMUqIdzFxX/+jjx8wRnFlqQb4RXQhV6xyG3M/t0p
BO4j9IowCWPI27YHObFXmzIEEwL9GfiIxiPc5mB+H255X90+fGNNiiN5G1U+CZD6
aR9QonB/3OqxjyR2t9TlMLdjz50Dz7Vv2Lxh68egA3X7LhiiMn1B7tysoHgVeRJs
V0EbzhlIwYhcQmfQtfKeowbVBMEdSi4ProPEdalChEpltIx2CD4Vs2JEZu9mUO8A
xWeRQLo+OIZ0ZhIK1ugm/gzkGJsJJkTtX0G9QZxtY2tdd8AUKT+7wpXDHY8HqaXg
/Ovu5ANsNieMn/jcUDm0VBIiH9J8KKhWjmmMTXWfHuOdfJh7NrlfZX7uKHV+3peC
DursUM/MEDGlmoG69JludBjLtRbDp6Tv6ezCSaBU/UAtDoIObqoixCY3JVL+Ez2I
xfRBxmtnsWmKFdwsu/T5DJ825UMIhTkI5hBDVvpvxXMR8yllA2WyPr2TbdsBCkPM
BQVIbXy8DZLC1/SR7Fu7ocRHbNrZzicXxKiWcvIc2jchx8DDphrsZ1JK5V111zTV
TrlLlT8Xm19ySD5fv3BhUED2tL/AQpSSbJt9UYCJ18pD/iFHGzQMoGIx24MT+rFM
WZVyC03W83Xbkpzc69vRd8IZMsHdQOncGfNap1WbbMQksYCBOXZg6jeMWNaF+ajw
imFr+UEOA5dTOMZVqlI8lHFddW7m7eguPwQjNvDLdp3I2RUBZFBsbkAo/wig1M1w
83xH8eTeSI+zkIrGg20jQl0idoHCaxSVxuPvqi8yF1JsEQxXSXheX6TqYK4HSowD
ZcmBAd8lboxVWxvkx0vf4hEMlvnB3xUZHVw1ZVIjI7Ne7X9TUt8zd3LQej0Bio8P
OBIdxdpAqKcROQbQvrKQiiZ5xZ8YWCKXNJKBiD61hFt25Hibk3qxlyDbFsl16Ba9
wMBn23fY9RARF2vezueW7K4c+Acu+e2EZHOowtILnOMltQUv+uu0Kp1pMx5QP/26
xVB0LX4akEW/EFRcNi4htscyyFcPZvIBEFMw5biV39cBsScdBq0UBPx4XLVFtP5m
qa+mb0mJRcaqjqKz5PNDihoSeCVIQpdw5NR23Am7jQzaJTGNm5Tu9JMR6PbGxCxZ
qazFGIs1fFasqUhQi9Q9oEJ61lToGIpk/nT6bN1Ip9fTpoxzrJpIUPQlHfhYfWKo
hUMdgvylRlZhi5rI+aKlXYwU/+X6nopdOTY8NzhmMwOoblx1VfZmEvVjUzILXfia
Zj/ppu3mUM3wkJS3Llo2uD6wx9cB2SkKkk0fbBffjKPuiCsXlAab9iNhQtm3Tl6b
AKT1HFZFFb/u1FmuQIY0HQ4VRFr9LPtgd+jSYfx3Ak/5iJsDj0rC2L2xDVkl/D77
pe90+a5/2tG3T4HUkyum0sllz+MbVo3f5rhii/DvOjNvK6+wDsZgr3GHkRXdRIWL
LTwzStZq0VNY8d+AW6qwUCXnOj4xfVVbbKf2T0zg4dFgFkrr3wEanZMLu+Kt1LHA
IJPOvrHwXUaZoMJBXBjbFpQSUcmSljyD27SeEGdT6v+Z8sFvILC/6Z/1BGwBzZkc
Tif0vE5dceCSGYUVNZ42I+Rv7ctiaHDJnTPZXMns2zKois2gw+B4O2n330yllzvU
1FmVzsxm9O93CThH3Ov22m2VNmDIZ3g6c1M+pPNi3JKQdhvTSlqV3+EmuBfnF0rT
nj+W5e6dnkrXMPBOUDA4JsAbbti7YxBOXOigly6ngx23IOj0jeOOOeaCKyyRYDc6
Bwtt66cPxzenj8pLhCT8RWyew6Jn3BBEwnfT8RKVlmyRvN7YI/NlH422LSBi7yuj
PNXMBz8V0lwvSxqxPZH/xeJucFkMZVCr6Ukx/FPE2nkEvTYf50Ab00kcozULd+xA
udRTNYLKdLk1srf+lv9ZABkhuGxuPwlPT//w1lDbW/cgBxbj3I5mOaeO/Z3wqzwI
5b3AofbwlHQkvTjjLW7obE5WSuByNyWY7PNZX6bSkaCYZMGf1J3/ufLB5U8q5BL/
e8X7f0x6EHYDdotRhoHUlsoMsL9EqJDPhjs8uC1eHSzlMGO69+2G3l7tXQy4YGut
VonteHZJU8uSDBMx/WM/ewuv+Uyj+xXah52/SI+EClTeMwZF5CaKXOrgVC+YK0MQ
clZA26oyX+4JHinifE68moywSIKtq+tZe33aTKVOfo7GzAV/yvvJiqu88pdTKAb6
f6iagBqS40QImvizD4T/ONEqXo52atzhz5VsL0ivY6KFTKqQhT2kUqwJSIEmnrap
CkAyUvi1/F9E234rm5/dkNrGYAigg4JEpbHgBicn39M=
`protect end_protected
