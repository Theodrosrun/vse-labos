`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KuZZr8JR3yPB68jSpiMkWiTA8rNzMagtn0a77hPJimi8RpZI34sTlZvt0DNZ7PsA
/qPZyu9vuV5eccav9JXs4j3rUF49TxWI550w1l+HMe6PNP+NBwiczH0bZD0hLxQd
INwgzBYpSrgSN/sj5X/0J+/lUT/w1rESoY1liNQuYEVzugzzjtaeYziKGDuy8W5P
FXJHPzcniB4o17+m6b74Sy66z4txq/JL3Lv5AmjzG6YvSH1pgvxsRAltkWlSfIuq
Jx85rcQuykQhWsdcs/afHBpV6QKOXWk7VpUm2SL2u3CQE7dXOrataEUPj5uUQw7X
uGSe+6v/KLfDcv7hANzY/w==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6368 )
`protect data_block
cS2Hohx7YoL3YmmmvhrITk+e5JaU+pSeUeSa38GqTQUlsZeW/Y2cFY5c2GOxEOxd
H+LBHOfYa3aPB4hd50rbVVO2TWKSXXKPANQ1BUlR0u9GnttaIrmDTfyQu4VlU/Md
HzqmjqfzYJoGsjGTU7bBQMx0bpQtCrKnP4bXtzXGIuM5hYumGEcDR5r2dQmWAYt4
uadFvfHb9ko67Dl2lXkTyCmIZQxK7xRoQqYufryZyLdtGHSNzgnBBDeEyO+pMNF8
+IGqGYbamQFrqWwE71TUN1DoSBf2MPQHTyTPkTzjDHMQynqAqVANL/42Sfxe9yoM
SvGS659CMB2HDKCmT5LwYRFpHm5DYvrPDPxdmykOKs1ONKS8BGCQZmlFM54zys1e
rlGvCP3bKKKZB4BXUbRv2T2CFtt+u0cT6LmxYFJqkvUxD4AvFOQfA04C2tYNXbun
e2EqpSqp1Q7Dn1Fcxpd7AbWLK9dvGzzhC0FkBx6hWttjN4Sr+gJ+fyqJQz5pE4h4
ER20fDkBiYorkak6jQftFNV3KM77YClKXhjperVpocB1KliHOuMrfcZOsqblHDs0
BVfYsl1qV58rdEKMvk+1Tm8l/BPHcSoWxMUCYyFRW2CW3rME4hfKEwCBfXz2daEG
z5SQutwTqmRHXuQY8I0OTN20kN6t5XVVmRVjw3ODr7RBbB1Ov0Cbq3pkauVomtCr
o5MHawHZCesIrPzOKJeB28mIQzB6RKneYwRtIHBa4vsvUWSdRfzbcA31C0hqSCo/
D0qruJQOPH4S3n4pw9S6vm17WnIrqqHtDACymzDK4bcXl3L/zXU8ZHjetLwlmQkQ
a2eFLU3ID7v/rr7mUbEPYUtC/njV11QkdXJ6/iOwMonl0Mnh7wIJT6Qo28CvkXsJ
z8QZNYxJurfo7vSd/qf61fWrKAFEe1jHVTsl3Eff54ZLG4/QdYLGvb/JEzxKgawe
GcHoRplXrPa9p2gQ71qgl4Vv4SqWnsKgKHtCdSLkd7KyOACL5ebBQ4AoEj1QI5rV
VLp89I9KHU1jnYR8xRfBowsi7rcbjwzZC/2s5BpjCHXgFaYX0SCXnQQTVBc1OTCF
Ys5HJcr1YFzMudQiFAlr39CRtDVGSLP/Q6TUBSTrrn9EEDYK/DhGIB5P/vcVgPDL
ywGXtJhc589YtuIUhVpj64dY7xYY+WWAf1K0rn9AXmtj0gPg8We5m0Gd5Qab2L/C
z/B7tCeeO5dFXd1QmHEP88V6S6mKLgcW+zXFnksmP9pnT+JcE8z/KuyEUBXEhyLL
UDPNIA7MR2OBXnrHgkRcQuluxlhOhGuwItGOz+C3rBoeJKem6rXG34i3VDZzTsYx
WwPZwMl/720YBatKUkwe6s7Qgg8w0sbSxLyrd6Rc6kcTIQJUvSgqxUOUKVPJW8PI
UG4zCTwMy0tZri0ZW7UlbIsx0mMtAi8Ox603gFAA9gVjAD21eYRmLUO8fK0OauC8
SsDe0nnGJ7XLBHnGWTlleh9S39XZML8C2aCJkV2xLra1SXsk5MhyZbULEmZWItOc
L24z8LyClEnsUJXaIqU0RppR0nhOzT4NZlrXLZnrDsjf4ein9pW/qD/0b7w2d/6F
Erlv58zcFjmglIEEW7BXcf4QIM/87cNW4hEcKwV7dXdgMr3zLZScbiu+o2aeB6q/
TnCURZHpIu6V1KBWPTCwmdJwqw70+MDZ/N+xZP8FS6w9jVA9wEFh8kl83MoIbwAl
jD9XFkrHNHUzjw15L4fuTgQEVi2ZKotzHFl9Zfd53RxUk4LPompRmrC6CeifdoFb
jisdYpD61sa/D/EXZZs4/G1QK99IeeLJTz9MDSCNnYO6vMtBM9OzKuu+vlqizHw1
DF4HQc5lnbiTZbA5F52+/WHPz9BIwLxS/uyB5bpxe9Azez0Ys1iumplN1HnT8z1a
KoBSLXbHeol+JsSBt3wmnOtL2WGxqPZM5rdlfs7gx+uJoDFPgrs20yMZMIA61Vqg
IuRej1qXyMu0jB6e6TwCvVlo5bUYHNnXs4ygnSTvyi8obdbjGyYj9vlVpt6R6Jeu
o4MR5Vg2xFkp2qaSfkcO0odWs+tP3iDAjAsgeEGtEqzvomsv0TzawuF+Qvo6G1wv
Jn/VWA9Tq8bf/xTi8SBlJSkh6q2/HcCJXpANhQlCMkDafAhsjk9G8eWx7x7rGcnK
lDn0z0ZVZu0Lotnpg9d0cLcULLbK1RxhXqO89dkWrAjP1xDHy0ADl+HjiIajbZ/n
2tLBvGNsXTwqb02WhVgNC3ux97hN3lk5kSLlDX6uV81aUYZXYqoTS0hTsNumSX2R
Gsxx6g6IuKLUMSvUg3bVSZOj7aqOWxEZD5rVNT1dmG0EEBN1v2HM2cPNnZ1qmpu6
lZUw9nl3Oje47cN/MntNT6o5EAUw5p6FK8WrtzdO7ojxJsAy5MH0M/X/mIHaqM1D
K35OzCARbT2iQihVDf/LWHs+AsGiFwEVfwv8Y11XfngsZ/0oIo+jfw335LpPmfpf
Yjpp3m3YbGeNNq3VBzfJTdIzKsIREzSQ0Vq/mnHBB9MBtrKScCED2LzQ1ZZomMkT
s3PowYgYh0IyzLlEZTWZTXIrKLgH5A/1ckSuM02Nk8s2v3GCPRUiS+67HtqOjzGt
0/TCDVutqkhBxKC1ywwdKUQ4rc2+6zU1qvw3icwwxs302X3FIDOx6Y3klaRnct+S
quSG0357jJH+qyYJnrnPQMZzq3NJUCzEy+O5dpOz04KUhPa7/y6ATRqKEU5c62hn
eo5jRQqp6ei2quVOGQbb2LBQjpM2xUM7k6gWr/UpXHZ81n9axrw0HF/G3xFOoqbZ
h814oIsxbzymkVwOg9w7gApYUaDHA4nJtQIIJvh9vZ//NK7ZUSmLQXu+aIbKMsE0
IJcJqGhUGZK+T6jW7S/xJf7MMIAJ6V/RfwY5s6hYXHglnusuqQCTnh/eDxQolkqr
TZy0UUT/42p7m72i17FHFTGg/IeMEv1YaDqKeQe8OWMyJHB/Fkj5QK7t9hxz7cON
pw7Kk8OJbPWsLwHuz0lgLwrv6Ue1NknG4DglzwTAO1+z2j7ZITjXqTYcO1mfcORC
l5fvn4EjMjOz80zvGqF2a0R7sbjPIPZx4p47a2/asnTQU0H+Dc/56TJCChcHIHme
56Eg+8342dAnAX8tRPv3/oR0anS80jOf1/jLHPudSFZgVI1ayb5J8cb2mes5IoIg
ZZfYCnqvy7/NayR5vhvoUKn2KmRyhDhkCbW9fEEWH/hX5V4RgpEfeJkI4Da/EdZZ
eo44Fb/CdxPADsDMXCEThAzS9zeNOGAWjqvgYoDJsdzAGZCbOnciHK94NGRJFktl
4TZ2O9dqYI5HgHy3mbLtj/PCn9RM3CfAwsMF61gxA5S8KvLbAZGTvwo0/J/nppRQ
cAxZglLa0ashxg6QCr3DXJqSqG4mgCCk9oTLF00h5j7JfFFi9rO+T61JCksP0U+v
BZvty4NqJ6LxO/xzFQj3FohiFXYgi/o7Na8qvM4Y1YoEsdEMylcI6jLPjWJa12yL
eL9thLByMZaY1k2A01E2m+DUOyTBYnVt1+9wDzJWt5C9m0+MFoI14L1b5EugubQx
awrAJuSZ8pReGlUiLfahfYknuznKBw2qIbZS78HiZXe3UYkgLUY660YB1RuU6rat
GJOBU6ou8vJw8XGuWQaSnp1WPRmdK/AWyslRMyvVzmocvc4a4dreyxnjSniEQgB2
jIFBPd3Cp56UO+olXXPwIslS7tLyUMBt0pwRml8j3DfC/IBgDBKFLJxW1ds/S7WH
SMpQrE9FBPIXkVDi4Yfi2+DrfFlUyQVt3CvO8QLBk+RNaPN/oT4kfX1jK4OTEmSK
eCWapfTYcm0XrXpBSn1hyyrLN+/HpeHkbEi0F2E89xsCgDBiYbl3ZvRgJbYXfXyi
fOhtIg6JVGbvg3x6qB+5mSXQMofZZnZJoWkheaxLuAQ3EHcUpYwye19blBf+uy5t
1XHrZmAKqLXH9X4+82HGO4ek/pfVJBAwfZf/bBKERQZDW24g3A5dzrMugdFDLUPf
i3wbJmvLWnBuUuY9xJtFd0qQo2gBzZuSS6yG4biXurH+2pcpJfrsTXeL1YZNuc5x
5ngLMQoJNBN00qFIBRTaFXIbgiY7WgKQxafP5VhNuW1S8xwqQBpAag1EtWIUSbvd
MH5Ga2r2eQleaH8fu6vN2+S2aaBcLeCkIFHv3wLwSyhEvPm/8s0iv9LN8D14YCvg
V4E82tG2JfLz/aI7i5R3e6osgR1/9wWeSbCo+HRgFj+9ib5vTZbzkreI3jJzqtMY
AwhBbKcrnNsTivJYxZsXBilBf7ZZvAj/0fMUVbxTO3N29VwePnzmP+mWXKwVvfaM
H/8ltWcgI+liSixSRStR37/o4+wECWAoShEt5fLDWk/sZD4nNyjevAZA6G6Q2NIL
uftIPyVpUmGz+NzQ+81RDVm7agIpD0Ewfv5pznxcB1Q3doROjl0WwJOxoCSgSJg0
CUAKziNINZ+pjaIRzNkWgdyu6QAurVZZSpNCvNVvLeN4UOgg3eybKWNMN3hO8G7p
Jrk2vN3/idTVL1MLxNnb48wCTz+Gft0m2fzWwmnOH/ZM+ik/xsmIsHX414CjL3C+
DjPQym7DCIBWl4KR3NRSwB5/c5fYgtwgIs38xwSOary0z9n3mJ8wzlIqMmMh0L0E
7OgBWvjQQ/QQ6MzgaKLs0+LXWszwVTfMipCz5exYaJo7fbGZ69EsJ+Tll+UWu5ih
ZIxjIfB4zEEdUPqYyT2UoRXp4+U7tdlqi7M+6XqBPfo3FR2VTirtHX7xK9oBKpyO
3fFuImlRACPZZvz7z/Nyq/sgFQFkVwQDnvAYZXi8FRvMfHAmZRfiTXLfVGnKL35U
TwfYVncxLybCiZRZa77j5JHpZeu+uMAkZMPgdspMoikjWEmwVYQWUm4fbELHtMFB
JEHhU0CNCA9RqX2JXptwTOB2ozqIduVSLoxaqenJPX5CYyvJaTzTpILyqZ1RYLy/
BS9EbS+stxsyXoklLQ2JjRfXg6EiPe27aetyFZXzMqO3eVVVxk8YlZ9vVVLsI0Mv
nfB5pHtUmow/tMFwF2ardHJEwDO0g+Jwcir7et4sY/4dCqaxhZVeikqkx56DtSPe
GKgl/UqYmPZlCmpkGptdKj5jEq5pnr1KZgDHcmsrxvjcsEpKLVX6fjQDqidfLrlB
jeCkZo4+C0tcrKrD7aAGIHHfe1MEaLxCrz15csIsd4YTxo7sTaw+FRGTL0lhd6pF
oHvBd6dg63NnuBB1i2j8Z49SsyTJJHbwomomBb1uarIDBNow0/7gCnQNchaW40Eo
o9rkq09Hz7IoqREKKMONXQyXQGbAIyHCFBwem37oTe4P6EUvYcYfJ7ujF03Tkeon
q6MW8QK+tZ/zgZquyg52LqEqG6qyRkIii0DpR/MLEPggOB78Ft14ZhNzzO8dKON7
zAolqG2XoP50PxUfBwHhafkQ5Ocs5paSlmOAaYCyUF2uiv1COZ8CAZ1IQYs7aZ7w
IHCKzeBbXfshV6zVZt2geYXXZL7h5D2Lgh2qmpnAi/+cESmQgz4cDQSKGg5+KUa/
tS3tsxa21/pIe9UYdgEkYjxfGuKxIipJqipVJMXZFUZbT3z/HnJRAlSdCqrcCV01
OLAJWSKvMrY7mvW87coqvmD/YiKrGGHoeNAeeSa+62R/bGGVLW5q/02ZQ84kw8zd
1TyOCyeaRzXYMG5zyv6tG+2jj5pdnXHtKkwh3ONSddbGqej4/wLpo4ucC90LUvpJ
gdd+S67BYuDwJgxYWqgBB0eBp09lH7dLfpORatovTtO3PH1xZLdM2zBZb4DInMBp
rMNgxdJAyxze7VamRWRmDExIDfHdexjVuELOPb65mvmRDsgzcPrCyoqIb0qV/CfA
V5c8zLDZREXYf181/fd91LPR+DHQ3wiVIDEGY9DqDAloM99FogKmDmLzY4yBUv3w
itaR3dQjOKPy/8ax+a6DAvjvHlDqTO8l16AZpMoA3f7wkSkbGz0Ur5ZlASiuQbLe
KozwwNdmIbBE3QSpwtZf6YR23cA3FmFgntTgLYsPM+VE9fpOXeIUr3Xs2YPwYoei
mqqamwAM+DHVsY6G5/KbuDGvWWrYxZNRk1UTMxx6hR+0p7aq93zoZV4adra4B/uG
2TYyeRF0IbJ1kwjwSWgYDI1l/nBLwpH3f4j5v7GnsTXS6cf1kOg1b5Pkb9ANq1Wl
61fScA2XANbcmaC4RRhiMFrL+P1uNb0uwYfxxdkNnE13gx2NQnpYfa3KfSNMO0Hb
ncxqyXlLjrAG9mAvh9vQ+lUuTRgTdWwkpChJxp47n8djWu7BuRzDVDinuZtKiHRl
ZTUTt+iwmQ79txozIYd2AaVhfaDsFH5y4bXt8Q/hZ0lYLIZX3sTQKu5qEMIOPRSH
zpiJhKK8Uxqy0zT8mXW/3Y35OsoI3QN3BYoQeCEef/TKev/ShG3B6L+1fmPgSTiq
HDPi77GiK4kPaUoeoW7r5+hht+r2W+5xhR71SuU2e1t9aH2q5p6Ta8pDEu3dLZab
IKBAiHOrGzZyaOVTJz2PCektpbb2m3j3H6c9gAARZF9ulOoPh64j7qaP4oMon5XW
3HkQlJtrxdCl4iN6YjfLBbHXcIRRomZGvNLOb/k7sCMebR57LZl39UKMExidQ/Oi
4gC8hgCndP+IBVC+mQY/NSnsV1CUDf2T3nE1/0ut6x3G+kgZpG3J2mKzAKIJgA9e
Xj+lS0f2jBT+Ta67E5eb8/FkGiMt3UE85vM2jjrLoGoHadrH2cjjM7fVJYpE5Pyz
jxH3fgOJaG8If6mHty1SewgzLc2V9yRwsYaguRb5pSe4zlii/AeEbe37slqnU341
FUZhe5Ta2wQ6zukOJb7kTO0jfkaWcrp9xJIlmOW/ux0DPMBO/NPAJ5cuPHEyNsFK
TjwO01UKN2mQ6oQwfowJSPAxcO9KPfCWmagDtQiv9UgBhCWWgyVGYImFvJw8KGPk
ZI7c3sjtOtu+C+oVLZnOqTsWgYHgRcFIp8j51McP/lvasaJ3YNlVHXt0l+0KehQH
E8KSqlURbUp4tLnOXRR8VekYcIueSfJ+sRO0fFNtAB3phoUmNsTdTd6WQ6a5706b
Y2uk+JUtiimX3Rn4+QrvVpQpauEkvaF+Ry21rnz4Q/Foafz0/UKfKFNa1+yizy49
yXydLEIFOjXkZFR7DN4vUgzZeTQ0kUVbioq2jWlacWfYi2+lGVZITvCCbg9n0vPe
F8+BqGLxKXId1CYRAbrEue9QsWAuJKjz31IWDnaamqGs+tdj/3mMOLwvLVkBQYgz
mXB1cbjYu19B7i7SRB4JRL3K/Cy9iR16cjm5KjaOgIeCVhaYAuVJHRu9RjHNperG
MF7zAGfNujV10Z43az7bSdeuzgGCE3BFoFgaxsRVbCF5RgnlmYDr/uPQxM3zDoTw
YvKdvZc8ROYo52bkg01RGpPcbhtThib78e5l4NpJ9zWYRl5FdNmD/qbrWu67KUrz
nnxu0LRVxfmgCoClLFvq4aMt0kYMVNsJ/g0A0w38UTiyE0eai0ijXzs2m9zKEJuT
2kBKEkhtmwXRnABnH7JKMnnEEdEyiNTOv6r7/MBBH5iBOWou7ox5RqJlWAmFTKiQ
iyGh7/ZTYzlUVEuFuEOTbITD330lKyUWJMTXlzKqG/CrHdpShFT+yjm+xQloCWrQ
ksd2YCud5GEbP0/85iu6N5Dq6UmVr+SQPHk6Z/KcGfTAIyZ3kr0PcE7tf5R+aRtD
ewTIcgS+I66pu9pB2u6wsnnRTSPBwSMGVyapE75+St4iazZwGdmbjnLDHndhlJsv
XV6eoytG+pBmDHlxnm7LzFAv+WKU2lPJkrqBd1PDbIyuW8ZdfEjksUML+tYyhBTe
EoPtJ5jgsBv3yV+/CurQhOneJSWHFav2Com7teM4Kd+HpY0jTIYVWqrMKpYWLQo2
z/H0m2K6Yu/x9eZItX5caqpEFC0RppkrAwWsabg9ZEOoX4vofSd+e2gKmgWH6p6I
x4bLqw9L/u8Fm2a5ZFAXuOhsY7LybzhElQVwlLnFZ68C0iyaL5aZciCABFYTr1Xj
U64MbNGk+ZcCXensfqGKwa8s8CGC9xHsa4Zxg6uUbCKs2Yt74P5L85fcq+pVH6AF
mzryEfM5/mwLbxDG0nKRBexEOl541Ki4WJ70VDW4uRrMi2XAdHKU3dU0jfaXeLd3
g0pTtTIZZuOTkQ5c7n19Uk6IhjdxXkZWmsBl2r39i/tnxaiO4dxIMDb3LHXPkxJR
x5krt3Iy/91CyrUlL61ud2pFe6gWICHSOwIzvly2ixEfXRDu3MK0ltr6LE1wHsUk
6sOfu5o1x5VoyGLN9untu1MtPfDnzlE7O7+4BgpheBuYFY5n0k/oZMzCfAz+hV6I
GAS62LLdAiZrBloDcaDs3CXPG2HNF+dRznM5UcuL0SaM644kflvt/9TlLuKYfY+C
gBv8/09GBZBThek+2LlZZyQjlImksPkSi7qlzEhNiMs=
`protect end_protected
