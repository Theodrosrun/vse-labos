`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
M4GzEvJQWF3MQ0knc06LSAiCjGcRtn7Ucv7c2BUZjqEjk1m+xFXjm2J1cxDQB8VD
KZ2mpkfZtRhe6st3Fk64hxY+iz3iv7cj2mQjWWs/I7bdxdcX9kG8atGMsLVYSsYj
alRSc03Nto/2w/He/iFDUtkKYmIJuu7e+LHfxtegBaULL0EfUBzCO1jtiJSevJPq
GbvvYEvaaX1dooL5PGX7Dw04hkfCW1kFm2jNXcY8awyP1/fNByWF9DmZ5G7EMK7v
mXQGmQQdZDYTspXFIEJgZTV72fgKgC8d1+1PizHb0rlk/Saa9RXYoLwVoXIorgNS
lBHfUILE1T3Wr32r6ICaag==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9552 )
`protect data_block
oiBvay/mA61FnS/zJkU4PPuA/mm5HdNPcGIV3oXEtSgkcg5lPTMtDDPD8p6sdjrT
MDBRBUyXgjxVqitgs3J2U1myw26snNSEzSlDm4DwxuU9SXZdjY5oyEwfDXluuTq7
WCaK1MKEp/r+btrdWxO0m3MQIX42tJQyZ/CDNQYmnMydenJ4eYMPV/Y8xPBIgVTg
FNl1vSAA97SG9v6fpQn1duxulWq1xdwKteIXgiRGGjifSH33c0KpSmCh50SWtjpF
Ty7RZXg6QB5qiA97F5u/v+3PFILCerPVqPr3kCnpt8AL8QBLQtPj2YWCtqkCwgC+
aKInkTYRMmIYEUfiO56HcFJWWjB02Ltt/TP8dSW11s4BDknsTIPRnXI/7eThE8sb
bsKKL8xBTcA9Kl7HqIz6ar3bajTpZdKufIyxvwSTJWsmk/DIPiQpxBL2td8tk5C3
d8uxaSwdF+x1wanKmAdSYVN6OtVRAO6+/s8xQGgBxPy/QFmN6zdkW5PkTwEgtfIH
WnjhffCd3lfuiguR2OQxeSey+4z8pegA3WEm1L7cPhopXAqc9RACEGYVuEdcXW8O
g6I3ysE3MjC5rnCEgnfv1TFhaURzJlhZVy5d1hxYxyS6LpwnGyzFfCrd+4hyg9ff
ITSpri2z4OGVOVWN+zoHHY7CadW1tJv/Usu5kyPuI4bS8/blrZXuEC1mlcKjH4As
416L7jb0vqhXyhX/Inkus55oipIiU6OUgdCz/O1UrpXfBa+wFTUtTgcLipFa5SWv
B3mQwIDYbdAjMx5B4gfZRjAXBbxytxMMLmKT6ehcbk2kssO4JJ+NElys/Dw/07dp
ChSGkAvlJt5OVESfrL+IGohGV3wtot/vzM3tIdMPTe3PVR0+QXT5K3eweNMNMMSv
TwRP+zJiTH6mNvIqmOOH0OG0G4vsVO13gXKXZ413uwbGN/9dQstrpUzqNqTDIawp
324O81im1uJSDy/GR0cfBwkBep5Iy4w208DKqx0Ymexu4uG3LaiJN3PoUsCdEw4W
F+1ieziVDBM+gazxuobf2EK6voKbupQbpw+nCRyrOKRHVlQbtT//RYoWa6RVffLf
Y4fWj5F3My5fkkM8FVlPrFEOcBUhi1zVB+M/9ntt3D1xtCsQ4Qf8aF12T0Jm2ksF
rAupS70uZWEwWy5/Yqe1qHvu0NM4pkQm5c0RfvWjcQZLsGv3OvWo78RFhgeALziw
nWIlZTcihXaMxhnrSQqPEePGKGU/yswrYtXL4wctUviLjH4aNs+pyUelbhwIyQ9Y
OVaiPg2cnsDU6VG+GkrJ00Y6Qsz3qiYWiNtxQSNWWfbeveRQL3gIpTsd+i/k6BTO
xZgvDDYN1sYTbvLoOFQ99+Qqvrx06BT3GHN2/gxal2gwqJF1PnbyAr8vSGqAhCgm
Zm2PcXdLvZHW8DmQ/NzmfUMqN0SsuUrsEaRnsPZ0OxvN9PZS4qF/bEpUYJoVtNZ8
jCZk3B+W1zuiKRIEQeVtmo+KZAJRmTJEfo+7pIIVigel5GUyg9JPKHELvvPCpv9C
jI+9yc+Dlufa/Uow3StJ/tNcHpEHirRFfD/vP8mN1zAxBxTlcrk2uAnchJdGgeK3
bXb/TgRLBQbk95trwWqBNdtuNv3bQhmX6/wayOzYKIxdv0kdyrw8wDkfFskev1AA
4NPqKCzZ8ynFFcndJf7OW3yumEJdRqG8OFBww0cPpooUJs3y/UzHoUnoiZj5Ak0v
4ANXB8J/Pi+4SNJufeR3m5tRVzwb8u/sfQara082/LT+CM05KOP/FNdCPPxb1Boo
FJ2bUT49T7ZUanrYBtASSjX39cduCqQkpyE8uVAugCC2sLQmR8iiqFMAJxfnpVtu
uaNnIXjgi435UoLNILRvgTUUS178OMWKAs35JlLWh8w/xPnbBKwN5/dW9gPlGKKS
AZVBKih53aY+PrBII+BdyHPqlfLBxpi+KIyZCqnSDmLopjDLKT7DfZxBXxWgqfeH
FjirQyLAdskE7DVIgUTQPUaRBBd+zVy5rJClwYE0JiFE5PDU76kFxR2PPXMG4MLV
VkSzIl2wSvfghce/fXamo7iYnYQasn64yrjE/p21JMWFr9wHunTg1gwA23Avtf3E
PHLBdYMlDx0Emm4rp+flvNeeGLNCL8++kH/MnpMow7wdWGdNxqVPyNRWanm0pCj8
3w5iJivQSBCOSDto29X4S6ZlqJ/yac8KZiQ8N3/0S3Ly0uk/Jgj5OOFK4CAA1kze
UMyQduZu93h/4X/D3rtVK4hs7639/cDPJVUFrUM308pPyvX98cJQN+ZvFADPhK64
G24WZRfJJNnJUJP6yF84jNEGbO6QQFLcoeKKT0gPQ9PVo+LhmeaEo25Yt/g+2COC
qJDLuu/7qrHxMX/1ALtCGFXriphSmdPvAPrVUdU2EfNgkbxOdBvirARkFiugGHj8
jv7Vy5ZSccyRd7n2zJSV5PLLD1OlTym3RS+Odn0yfpJ17dLGvwR2PTb0jDAvN4aT
7/ia7eOzHoEhe+f18g4RIeYofyeKEvCWf/w59fRISAjnSCFb57jEA+aYnmU3TtPw
arIWC9av4YIrCFWM32RtGWMDQGixPY+HfU+80oArNdjc/ftt2nTkjb00PYEJE5PX
WvSfSX+cKpOWJ6vV/3h71jTQpWMlInRkF0C9pWNYU3q7j4YFeHswPAcpxvts963L
wahZo+cODQcw6vOsfrrVtlcDSx5lTncw6xpily0AHBzt665ced4n9DCDUH2/FXLE
8076hqTfsccb8wYXP6LasC7ogTDtYgjp5N49vj9yGvBRspawHc9d7snFjDem/05i
j+EvFeN28+7z2XcWJg/uqS2J4NkUcfdRgaPp8forcpx12FhEaqnHBePYlSBduqD1
hkOW4C2JmgSUZ7nas/DSq8nFr+ViXOwvgezQW9HeERwzgUSY16s8m3ZX1TCWQtUM
UiO13sgDkbJ8OsDaE3XTPgGDO0EBOP1BRcjquD782/PR/K96t7v4uTIAD1S0CakB
wARUKc9vTH8YcHFm+kh+OM5tuQ0FD5Z8DZD3OFKfIQBw7LqnBaHJWtQ8QgJ2ZcrA
M5oNiSkj6GmYDOnPl4XI5S138DLMsixJePRFwUqVns06SbUFMWWUk57UPdfrtRat
ujYPBOpnxSQvhA9gP+EgLPycACuxC8jzntCRqy5BN5eyaMHGaBeqIUnCGdo/ZLDU
hDhuRZGpsGoTfTWkplkzwZj9tD5Z6Z9NCw9xfCRTpIi4X82ZBRQbe9DPTEb/fGNo
BkWLyxK90QPZVmPxgVnpcgl1HZWhCXQEqyuF8OniF5sYaoFUcUVpgChRsgap3gtI
jz+d2n4G/iy2nF5smrxC4n6VcejxKw4yHlyKl1sB4kdNTG3logYi1R7zqcD+peJQ
iXDxO2Q2umelYrApocgIgtt5ZTKyAzJxC57l+eyziAmzM+PcaKUlCI5JHDmtAbQZ
JOb/Y/AZMmraR8NHdCHM8BXZewZpsTAbXxtbf1ERIvJO86rY/4UNNkQjJfRuT7Xq
ravJzl93I3wMAXEVoYvYI/Alm4tOcHnDjzM+LaKyGzqbuWwEYARZAu1FT1TFGmYR
hLWoWrdqHMu/SHXrY2Zqyn8EGJmW7wkhfK7mbf3MN7T1sknXYAkgTdRkHM9RY4Lz
gFLtVtlGy19jpC48NgLEO3yNC3IcXRXZ35d+gjrht6vpEpMr0+jce1DY7mLg5kTj
2M2weX2EKX8Hhp9d4I+7XdnxWTLYSGs4ZxgpT1E2YB0pxWDI1l6rdPHxoj2Y3/7q
HXCeDlZPVxI5NycEitKMf4PingdvKg83Rihne80xdmy0xlH5XAmIJH4k5lLjQnNJ
ZMAalh7epdSkk3DEbRWfbrTTj90rsoIGpeN3uZmR99K6/1pv6MGiXRiR2t19e0O1
EtV2f04LpFKQh4EwtSBK5bFp6s00axcDwuJ0Cx7nlzJ2WjGhlmbfWXS+W64kyFHI
Dg8zEIXRV+u9daqb/UTag81G5Y1lJeyPPfKp1r98ArAUNRzJXquD9c9XK1iFWtwB
jiYxQTSSNhHkYFHgbyy0+xMDtgsqETVDltNoZ9aS5a4ZPQs5F7KPV/EN+3okmQG0
tfQb4XfpE+vKuNdmF2T3w22pKnLWAyDAvztKguyq5jKlkY6UmEZZCk9DSmqhi8rz
DhCZW4jEDriDbHg/BxSanUxkT4YKrvMEdvoei6E4wyqF7a9e5/kgLIVDY6vCUpfA
dcgxw5q5cboUqGK7/qb8X6t6bTn4dU+2aC9ti93YRh3tTA8JZnQ9rssxTjovoLu0
yK81/P2nz2El88aSB4pnJCI4Z2/T83GjbC39OC/VB7HpoQbaSM2sB71V33KD9XAd
cveTdoVxftooMaE5RxRqvjRkELohVG5NPb4g2UQ1ZGnGMJzre6RbYeXdVpe/VTvj
dTkjfuGcG1C+P//w6smbrphBOs4mBFffZ9fK5at6Erj8+regetzFpS7WlyVSbnXN
lQaf/VIwxmBEnNVOGBIK1ds5GkqDGoyw5uzlw4FyZYgOn56i2arRZWd/qSZHJ8iY
jTovPkZjze32DO90WSPWc5TAiFjqJ5HpshslcCF/RH9gXy7S1eVyh6dc2dAwg6Jw
ND/UImAA2NVkCxnUEvTJnzsnY9kGEYHSNDE8a+qCNjF8obbtNdlEmeIoY706MCi1
MJDKZMU/BGzjUMZPg8O4sKP7k7F99A/WV4Edq++IZCNycPrWJ8kb1IBTo3+OKa0s
7Ki72OxoUPuF/fxADqvJD00zlBb7CXD4LEd71OdPKxBZAfLyEEMbl3k7hWfonfJj
s+VxL7NxTzxaK+/yJbOIZfgGQMYuzcKVV3WDcN+t/TXAMkBwfqq2dafCVBVUHz5k
JpK5BbDs2ditakKby8A9SrDXwXXek7y0A79wq6XCKRzt2H9zFJFm5V2tlHb1qoqo
V+hoz4NxZs3mNx9XU4dPyHjdSc/bqQd9Hdkgju7s6se060N5wi9yTmcfQCHRHK+7
mn+3xRZW8IzbcED7WTYH2+LFEfEqwCFHU7m19WE2SBQhS1A6CqUxBpmhhoOi7SVk
ba9f0syVLb1YP1ITzbVcTfiA5idu667LMbRArDZpwCZ4RgE6cPBd8TkGEB0zuEeA
3MPEkj9/9ISIOKUIU7zMXoEbdSwon2WpagZZjK8h+rLk/9/nbRqAlcSOKYPLkNnA
m4BT61O2SlMsU9LcyiqL8k8I22cWWFm493lDtjAJUG0r9BLma8cUHyp8I9gFNZv0
tM66LiWAgZULWLEPlV2gdf5CVHoFfE33zY7w8IdJnNxN2RwFdS2YFzzEDHreSQUB
agMy02JSaJEPPM/3fyjEkvXsbTkDvzyRKpgW662++UmDRo1aGMeGpCTgMp+Sz/7O
5d2Roh5nbSykNUV78gzbJehz3FPfv7hfX8K9uaNjZEaV3lv4N96JKbbyeT6iLwCA
6IiFcHfG5tanINnB+kYVe7z8YkUXM5KDG4QHN5XqwwHkincTXC8dKJLbvlBgr07x
HXt/dz6xF9RnWhp2yGg6E8qzJ308RGIbyPWAAqmih9V0PrwrW0XwU3czeaxafjiJ
khlh+rAstozeC+NvvOJTPrvTyM7ZHuQz7mzO5U69hsUhU/gPIrHqsxFbvWI7fMpB
QOgRtzIlXQyfElTGUgFi/GUX9pqiuP2xW4exELV3leQxcmBrCqYROqMN7urjGtgH
qrgvK17vHUvVj4Lhz7BJVm+nw78g3t7Lgi4CQQGIhCQCYXZA/bLF869fPpkUUteL
gqY8rkQAvXbeJiUdLN1R0BvNvfTZST6crUVHrguAGUMIgdDTYSexBRAPuUkXDmvL
LgAzkircTxpqJCb7ZA5nOe8XS/W+KLZrE6SiZHBZKqaaBMAIwHml634ZtWewVnrg
JVKeHvlkeJw0juUgC2+cv953sECD4yQ1pbooiUcg/Vok8u7R9f6KpOgdPc2MS+wc
P3n7KygDh3PurmXVed/OObuuzwX2LBKKTU5RLrbdir9XEKOQMsmg6xVVpRU/AROK
JkU7gYSy9jHO/kk0QK/Qi5xB9hr5Qubh7KgjnZxJRppaI5RWanmRzXRMiLlfjLiM
9FdODctRwtO+aiMEQS9TuweglqI3GDN2NrEnAXnq2QHREq47k6mb8o7iYBESLUKo
ap7RomlG5QgKYHdkziTWmmw/dXnmDr5C66zLriZT4xyIsdAzoKtnGzfP2m613wg8
gAZft3AxLUfd2TfFJuBgdETeAq1KDeI1xXMtOg8LDhTGeBpMM0VDZeJ1umw6ea34
yCCNGmW0K2YEzPGxx7EG4uAvF/hC+Sh3nelDa9/gCsUp/9YGi1e01HLoJaeLCtpf
Y5BWblPmzWNF3/RUFePID23Mrnq1KwebtroDxoNExx39ufgw3GZ4zFsp+FCV7x2r
fTJXNLgFnApT9daWOIFsDBXwM4NDnTOt7AmbI9Q2uCCIEhhLRGPnZJejcmIYmtIz
4JVxbME8qCIwe2LO3y01IOwMgksQDxBtZfzbwhOn3/lO5zCuRptxnWtAQDRC+Dds
v7Wdk+F9KaQsUQeZ9MR1ieEMjZgezuzhyzQwK3thr6XRPzUOg8SeAvhOKuZoegH0
ASIVV2hfaIAy0iATOZNmJb7aJeC8a1DfXFWFK++fm1MBPgvT+ZgJD+2atUBdhsDr
L7f1AmFkjudvEFvyuzL4tySY542dR8bbHo/Kv5XI0P7sWuIpo5s162lbylrFTPlp
D66hvYTGlzvoKLJDmpI+PCldyprpFV1/P9rLjdTn995dsrjxi84T7VCGMQmbZd97
4J/nDNeWu8zQpXKfNZr73q778hXs7DzwMbtN4wf4zcpWBqUisVRn4VnDbBXL/z4X
r7Aodd25vpYF8oLiQoFcGsy8XfVc5nzbmysZmm/XneApDC0EauVXv0MQznjZgre2
WgO5j9vAZdBx+GrCHn6Fllj7wTgaiECz43F1pjDZF4rTF7g4UDPNqtTmK7s8ojvs
s6FB1N9aQdq6OgGxG6ajQGCc+uQ//DTCy1ClWwTSXtVg5B6RKwB/J3GeMgqYlFgI
HCq9Ym1gI+6vb35kOzjd2tXoLSKs02bKi3nfnNmmSkWC/dHe345nStYoVZKr+Ke5
Ptc9SoSMod355ySzxf7DjgVReZBTuAZ5+A7zt3JhjTyccUFpn2XmPxlKeaLCxz14
lQHEFwgigarWCsFbLMqFF9Y3PDjn5pTpqQg8VJ5vcgtG5uN6OBYVu66x8stZoJxn
QECY8Umo9ddj7oMqVwD01bIuD50d2iE6wgtb2LBE8yXmgcXwR6xSDQtBiCrij7aI
P2PwvhRsBXS3ZbrI6i0VUzdStIoWhv+fZBCd/oFZa6sBWwC79fPRx9a+UpwT3u5a
GJcKnIePFPJgRdXi43avquaNOyI+1AsuaIOQQAzNLLiyDL3nq0ZIQsWgD+/jgs5C
ESBsrURyOIad/elDapTeWaLLGu5tZucJWOCu/QJ3EkTv/NiKRND/KCQa54ejttmT
LKsd63rtSndJODEx7UkKBy5vbA7KNhbWSCkYkZVmRBjlx4x5FbIfFPX6XIKfcDgZ
iGYyjxDMix7mk0+Lq1lUxHNA1//EINHzCSIWu8vDLHZ7ydyirN5ts02HdentGxak
lZoZi6JEv+5DmYKz2POm/Bcyp/s8wJWHaYIRukGpL06S81VJhZGxsz6LYMjAtlns
AUJptCQy4jg1Ha3uPmFWZQqOTuth9bPMNkzN3zJZq59LyKsPUrqNjw/3ITJc/Ki5
8nc087/driRnC8+LOylwofSJfVFDyPvC6w7+jpw3/CfftIlcY07+hZQj8U5khiRY
QG7Q6Ik2aP1rqKZftbU0JRC5zUCuCq1yZkt8/KB7uwUmF8rTIteHdBgh3bDg5D/3
gp6/5zoFNenbH7rZXaq5TpZNZl27JkLwN7c+BempdChb+JmSiVtBBBBqbvn0K3YG
gklc7dTP1RcKt/NhDfinR9iGng2pn30WzmSXser1Pyyrr+ui8c9+MC6qeRWtRMI9
qkua02Ne2uYQCl0B/muFWQnBdb7TcVFRB7R/ZAn0O8Yml+JdvcJMlubQ8xIs1EMW
Ld1D3a9IhMiQ5tKSQU+0YqMZH4ZLobAHsXMr6MVQjKgqcmu9ImtUg58RL2IdbOkU
vFOj/Qvj3B6X4rGlr7nq8vxsCBm2LP2B2CZJuLiuV6KdZNvIWz4IQZUWgi+uy4+v
IuHrgF7iutswy3lnZlEveGhpecfDnHkTmGsKF+ARRK36AV5NgLCdP0HJhHqyUUwE
PC9gguRIUtDBE64odjLENb9xZH58GEFP3jdgH1RMmVXKPQlSFoJZTyUMQ6W/SgxD
WGOaUja33j962IN0I3Mzl/ZNl0mkg9wvCPhXIR7LndmAOpPzivovFiH21WD2yx0j
+ETeUuNAAsdX1t0dZKq9BH9Tp6VMUkbtVW+Y6aLUybYyyPRixhIEhl27aU3zCTdn
tVJjZqBNrK2dBlVmMZo8b05xbHYHLb6wIjS2cXKJYaPVfVT9zgEviildyYfRHp/X
AJ8u+kQbAdcBetnnyqq8KRrtLWXQgHyOtqFVUbfvIJJ3pXbiJu+q1JBJSJ0mdnED
ZqsjW2IIhCnqIwoa1oD+B47S7AE1KirAsYGqOWuC25CX0xPYo2wOqidTpSQuzlT3
dNrHN3AN3rcrJZRxuPmrjajSh20kjanU0C6CtuXLaVMfdHMpLTNDOUUVealZ7gEQ
APmw2hPNoIAp6KzR8NI2CSPe1U1ohdUfF2pS8e7Hjtd1bpCPvfOOpSn68DeCc/PF
Us+uier8VbeP7vEUzZzN/Bi/Xu0G1mNGW+rrRMZeFjCpXPSjl8Sh5FlurvSaTQXZ
bpbZqSqMXcWCSSACCxz1U9S+9X9FBiH/1bDMSiLf88S+heqk5LwUCs5n/zjXrEMx
7KmX/NDpcgu+HdGkzFdDdtljCauYNr7dYhMBvUSF/aTHEKUky74+2OJXnSsmXyOo
+upmTJsTiRSTADCPwTdik1Q8SAsYfBbM+GbJFGIgdt/hYxO6fa/Al141oWEqJtX4
BN7GM+Yt9hhYfj4A/MR8jfmSAsAHbcprpjBLlCt9bDd2KnG+570W5YrS8myYi9IY
BinKmij4bj0Bq7FIMoAKQvQpvk1A/FVgWXl3ZP1Yb7ze0Dad51G9ZRja7n3dz6aD
NAByG19DNlRdQoS/Aqbtephh/K9s9WJYHHrv+Mu+q4Tr/tlwHG1szajR0ZTG2x+A
gK3fIL4vuqNtgAcnhMUFYQYuKOWxGSgAnToGxDw9WW2DEFe2V07/8+mdPNbWMfWO
lAgExlGcfa73QTntxIo+bg0sAJknuP0DRPw5tsKLyLUj6nr7krM7eHJ2eZMyGoVI
zUAR2c27Znn5BvBJVQRykDVf5zh6PaUhLSDOqK0RfKHFKe3eV3IwCjfQcIfhCHrz
qR3/i3YqxkzMrSpxDXapKsNq5xL882uSzc9ySMYvCwdCl9TTjMuKMVdA9gVw9dQU
fjNj47Iv/9LJSgAuxOn8agUymqUIIocaW3/r6YQlPhrTOVr9fH6h8BR6NhTusngx
AeQ/Dsx752LsNshzMM+paHUwa/rcmLrpE5xr6NfJy7BuldXnxzkNFcvjOfVkC7zW
4jm/JC6AFZN/R+jxkOUxQIHXMyU3kpWxkERpNBZQanCFnGJO8EFq9QgXZuPU3RpS
k+Y7fdjJTYZz6jr5iHQnb1IvBZfP8hL4m3Wjbm9/Y7M6/aQA6C6nNJI3UYzmS2LO
TXjqWpqvUbzfgefG6AnDLbWFRPLHRKj/EN9MmsNxpCld79QiDHte3YADjG4ydzWu
sZoQkvrCpbGZ/e7IQslAzxQ3w4DNt6YPRsNZ0jM6wZcLWDZSTsHzi2O1Yg9sP33h
mAzVczDKyeuhErS9rXYuvCvBwyAnLYbN/e0XujuqFybWZ4mF7m/d3j4hklDCWx5f
MC16VcsrBaj8BPwIofjR4fkNJtTaYyPckuMBYu0LtalUSisixCSEI5iUjPfpRQXv
8MzefaUrV1Jsc7jp+twwcw2bF0JajLQIV8iuMK9nKzm/2X6eroK8BcjJ0K1xd6yL
dFYr7AF9VYwolNr5PRvA0TOD8SD/kKSh5qLsWqD74KM0WbD8y4T7HOurxn6XJIlj
6kwco5dqmfv5wAt13Tbn+5k/bUtpDbE+ykk5zqhOAOfVyAmsnKhN+ZuDzbFWqv4u
WZRsMe03w9I/ngAChYbdsnDNnm8dxrKVmIzv9//UtiFyuVUa0KIsDIfCZsDF5EZ2
+MKKMzWMfnvw6NoseOXxjqL1CyqzDDUnYqVtN5TD6nFrPGLHKoQnOWJzRrZSibjb
Cfv8bSGWzon0rhNWvqc3O0m0fkFgZb4eEt7Owo84VSToEPb+SR9+4lXkyOcvIncu
RTtq4nimIo3Xo8hr0w1NxHCHINlgQBgpndvZfytYbftydDX3Qs1Hw9XxgT4nE8JY
ZaaIM9yC3/OkHialCseUrJ1bAkHv4LH42yjzySanb5fxA5THhwPP+c+nPxDCHqRe
ABhPsBI1APNIsr1ElWjLTbn1C/bptFmfgtZ7+sZr9i3RcwZOs2IzYM9/zTrgwiwU
qrix8qGwtd+/MwUZOGuCxKCSOFRMmptwn677vbskxYNXv2OGEmE3kmzQ2lB4JKfd
EE0PtQTNlXx4Sc1LCxNhsuGZeATsMF3oO0QgTK/4xiWs68XisDASZmBn3VmhPZ0B
1og4kKE2DBRG8BPoxJKijPOJtFen3hO48UQQHoQic9Qdhyhao6NOtN8Qk3KBCgA3
NUVa14UD+qKfcIYQh2l002hKpoxn40vIBy7wUMJQqhSL8kAcJP3uW7lCT8ZhWf0g
xXYPsTNylfiESV2EyK0lZbnxj3m6JwQBfzd9sDVcrOIzjmsHScGqgZgt/41BVP0g
bp+SrliHF5utrbW2hOfLe9KusYKIslsscKZp/cUAuSg7NwYOEEf3k9RJKeA1+5IA
AiWBE+PXLX5Ck34n8fPnibPt6JOf+xb4K0UtJIYvf4GOQs/d1w41eGLDPrmZiB0A
ibwQyoWDwxHlsemwsbFicKkYOqoFehm1KfQh+Hzkl9jyToNYSpqEhdo8tMoLvaSy
fEmTeTwrMb4QJySFdD4YweayA7Ku6TqjTGjtW99WTvs59DBxFhEBVWqKQolCAo5U
klLJ7y47h89RFUIbzFIgxRj0M2QcUAc5khrsx6o1+C+ls5gKwNyM08HqyZDVoP/l
dm3LdxD1jWHlXD5n3ux2D8Jjo+yG5I58tbvGQnh3Yl6Chlst1wONDHfVEcwiEvND
xMKzLrBHspNcAK2Z1PhrKte4P5SayZgKJTPlM/TOZbde2YtlbB72MT0g4nROSVOz
AnAZXzq/kcW2cTfpJPjyQqsFik3lSMpqlpct1KU0MWG/e4646lfCprKu6bfHfVfd
oulf+iGOuq6I3GoiDai9p0UIPhJM5abo58sTw1bzIzvT+GnpgSON8AgK/dhKGizT
KZDBLMrelbdhkHXgn5ZmSJFxD5jSio4DBT/pePH4c0iGFyzWhZmW+KX1LL/T1H7w
ssZXm6jMgwrFx7LovcQczeOawuaqiB7yJ7HFtmzpSjy7sKoZW0YJChQ9qLPU21M3
sU4WhS//LKGUzOxXlDrA7yUmKAaYDA/HCBnMPcwShYZ3sTZmh+KDkSvIl6F/kMSq
RrMF4BtHkybVFKy9N1kYsd/yRoRmbX9z9ub5a8KnSugOJ8e3eu3cAtfjO9SP0HrY
JcX1J7sB/da1q7QqUgSYP+1VlEroCYmHWWxNKMcl5SmxAY+XjD48ZdOqCSeWfnI6
dBXbEyehxhi+kiIVvzq314Uw3TGFhxzeS6/bpNsfbMruDV2gfMODOjRlRbPL6/Qj
pgPBHC1NaTzCl81IbGJ5jw05c58XNw3fGIEvBdSWCt1ZAsbKQDr8dQVvxaX8qHN1
Cq663/Zp5jwtLaji7cVTad0RT2+W7CUFfXmxQUjWj1Zz46ZQe4k28lnWXa3aoTFj
xtVBWfOrRo54zAbBOSjwe339jxJTdlBkWYnesjX5ODkrx2BXBnFq1hsCSE/jyQXJ
Tmete4aA/FeBLEWSpnJ/kbuFinvx3Csi/iUcAg0OpvE1k7d17nQ/6YXz6EKLwsLC
XdhUy3GgOny2wt056mo2uVmRP0VjN2oDDLC0w9ipk8nnRW7lAzMnXp0+0nqxGTJq
li2QNNmWgDZf0YTkwsi4L2VbsbWqJd1ieg9zTyWaR4FSOCcCn5GRDko5JJ9lWmao
g2RCm3MpdMC4Nfzd045oBit8jC1quOBJVeJvHaL1i2wcrgOZYhdjcTPCw4QN7UR4
6cwnlQlllJEB3hQDr3p9axPeGgE6ESAs9OD3slP/ucyy4Yy0B1FFrIl0tSBpfBHz
CNIFpMstyXG8V1NvEXUZY7mP62IOuNPDrClX9HYRNNXKDtnRfvo7sUGwGawo/bTK
5429GIhY5Xbg2KShZ7fyeKA+UWpS/MS2bEiJ8IPOi6QVqt89AJk0sYswyPcFjR3o
skDubS78CkkCNIr+jx81Hj9968qteMZiFZJNGlg+JbOBLzFhanYbr5EZ3jXbkLoa
27s+dbhjuMbbR34MfP7TYqUuPp+HXeU7v4WvrmwSLCzHmkcRVozTx0u4YN2Xmsyh
pYSI/FkJZilNocqwlzp8ek259CTarsG+MQN0SUzB6teY26HxiP87VHzFlJQQnWQ8
wt441eneCIf3PXgOWFSxq1xPpvf8U9RUh0bDFZFvxEHnTQ9qSzyNIO2TagEZSkCi
`protect end_protected
