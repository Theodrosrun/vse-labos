`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
nu2hUiHCY6y867QkDJbR2iZVKVUy2wY+7QiPjgqP5Xi75R2q/VUWkM/r5GIXKmzn
Iilscvs+IPip/NFcf5GwYsFUdA7jCz/audDHWxLA4yKunKEt/R/DkTL22p2V+BqM
WJlGlweqr4luE8m12wbnIK63Ies+PptvJ2I0VqYbJb2xelwpNwM1lVZWr2ao9nxn
EWBH1iICeSeQJuMWa9MlSpBj6wILwZN5rM+cKbdiy7/zMPDq9onjz40MVo3p+Rk4
ii633cjl7DetSmOt/05DWwaC0HEgx5XE6zCCXxfEvFqGRcAjA+czuium7kGrw2F3
cik2pV9XAhLY/7Z9qMjqnA==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 23568 )
`protect data_block
ihOQjCWx1cWbhn8hH9QoWRMp7jUjFzWwcMUvRPojeqVylFIqK8G27990ifo9zCdK
jrnFP7Ji0hedHLQSDcnVVBmwI/Yiajj3xhGsYh3aDN6JgQHJLuHwLyrZMqclOQ9R
IxltSoGWCPqyNKIkcWbM2Ej41aagzZeU0nAG7YNyyHKqDhz1xzVjgaGbJY2bs2Eq
2SF5i+3lTsEkffiZC/wLuR7P09ZJcPKA016ZLsshoB71D9ub95hzoIzlfuX3EE/C
1Xyf1NlUDTzs57OX/AoKeF3noGvXvMa9d0FqulDzrt1W6jcMEOPGF/tR1zFtHWx7
vHg/lG9d/tDcQSfKtjCqzBnC2rPvK0j0euxaGSlbAQWy4Ww4fwSyO/6nmwv7BRRS
7PyW/yb41Z6rLDBWdUOOG4OUdflLSnEgEi8Q04+WsF8i5f5xU2M5rvn7cEmDbYyb
AOmCs4ODre3/KGU4MbDMiHDxi0Dkr4kegXIYe5HFem1cmrxxEcvIFKcZqp+x7k1u
HPwk6Jdjoq6Fim0jDK2V2t9zjw79QLlL4WahKKhRpGQIXX6nMWP74gmAsgsQBE4J
1mb6/1q2IDrPquaWSumq2RnxljtQXf1b+ovH2iEWdCQkmoldeJ+FKevWPnvvkf2G
l9yic1HMj9ek26MhKviC7Ejj/u/eKowk+Y7eNYG9VCG/5sXrTb8C1a6RpZk98UzB
/cNoPnpwNwg+TfqDkhio6YXN05Y+VyiExoMa/xOUvNtNlNmLSxeqEiaHY9UnDCtc
wMZG9NI4hPjBUoP5FvoSenq9FUU2SL+GwAH05+pPns+YzAybPDkFHJR7gCnpJpZr
i/6hCkxQy530/on003i2upikCJ7DbWB7PuCytH3CnqfhGvtfDKdMPMKOAv1pQauS
leqfkHTmcUJZbBhfhQTotzVIMxz3n5TZciBG9tbWbZDHJME+DS7km3MNKZMkATT0
J3H7Ui2viXkLkCCDsAqAlIdTIAKy8wq/YLPGpErDiFA3CnB0UyxR24L2liDlYlkr
Kvhk15w5Rz7IOWZJxoo9tu2hKDvgt5BYOXnlCwNdr92bqeQlQsJkMM+dpXyGRDwk
ejE9BbTDdpEXg85A9HDUeIr5s/eIcijGVxxD51eUROQSjfeFCX3o+0UGo5EptrKI
mnghfey6zeFAYrHfuQ9V4t7r7wnXswZONXLkcH9OtReRUXfGEIoIkEW2g3fnuFLg
KSc38DvjVcm8kkuUBOF2Xkp0aKLKrhwANC5u/fB98L50wl0cqixxvwaazUBMBu9w
kSFJ+M8PVdFOmGGdlB1k7OmwQGXDOOMTuiKJYWiPSCS6s6y2IWqm9pl1+NM8TU0b
MsfdHZUHoWuNuKP8vqzAcQvaZnnqy5KhJh1OqfyUhzWd2blJjHMprDmjRcyu97LV
7gbntoVWTU8T0PzvXezptYtLrSf41acqQRqgnP60j1DWemobG7VAoEyAOLFiurud
jKVWyjpL8M68gtj0QUzKsH59E7iFNPF99FEHCWJpaDi6WFHl+jSczUB31U9iyt1A
kHy8zxCveldxjINpCL0Jef5PT8q7XUcB6GW1QpoVlR2BlQoj+eGSGnEqjqHuwKlc
4HJaIPxWv23eWQibVmOHPzM07VjwaiV/VOpB6Sd3k58bqbaJvNXsrxo4GVXktpnw
WihDnA4v5AesFLFkfr1aGuJK1QIQRp9jG1VvjtYWveRf22vCTmHXQCYVueVWSKWp
wJ1bQLco4MsPwuaovWaiD5gGRh0d0L9sSCUdOpxhnMYW24iASkBF6PtlHAU0UsZi
1fMce79DKEcGrqHn7OtxnOkQAuAAYknih+1PWSaJycvH/BoXeET6MbETdvnpwfYd
T1dKWC4EapMmzRApC1mFgb6Lvqz1yPwYHFIFpAdWDpfQfPhQNBRzorjrGKyWeAol
yrXs7ZQY8bji8hepXW/REiOS1mneQ8VDmfwNqZOQzhBuxEUH+Lu+nHOHssCU9d8x
SNdoSdzXCBDHR40lhtzon0sY37AJa/mBCAKg6zWWjf/ZOWtPE620wCW4uKL0qVRT
A5afEbhFKa6YKVz3txITe6Q2PuFfFCR6/g/AhjwNeKcAn72ooFByefhjMUkO2wZ6
dxTQBrofX62iEjYQsCxOmCIVG3mSsCqbncA/hIZFqxB2436CWLbFE2T1X6pT1zSV
RQfq6aNKXzSfheQQzeNSPCZfbN7l19HA/qcwVC6J4k3XT0a68O2z4hPYEbBAnjCj
NIXp9OUVCfDMmtBQZY55Rw+qpp5v/rdahRgbdL7o1ARY1fiapLSsNzErQt8yf1uF
vmGedrDoPXcSTgSoWdwBdPLKXAZqpU8LFUoNfDjtOKOhXAk3hEA+K9TDOVqrHfUa
uJy/+1qD50533gEE0oxOT/HakRdWEO3trsOid3A1pRNTo6CEmjPlDvpSF1RiwaRW
2wWPGvl6Hidw8wndrMoziwmxLl5mwXvzqYVQ95etwGhGCQq7XCptINu88u64sB9U
SFud0CHYiK06nycTg3MER/2yjBVmfNu8k4bj+X64W002UZAQqkBaOVySpkCfSe4B
PVHFWfKejhXlTHxX+Pqx9YlfX0s1Jd9JyAmXTCnvHV0bsGCg/5DiEr6V+t0qcL+Y
4Y8vhlPwbpYXIjexMU1rSSUJXOXypbkbIxKgCpYhU27GiqzNXHzMk9QIvB2HESOM
B0I0i49bL/70nnAvISvZDlKEJVkceRLXKu86jRzg9iysnOxefquugrvHckTgnWgN
jmcqgX2Sg9h6zuByjLZJzxhnr4C+uesIs4SddHjdgmtQjWxS0WNkyvBRS4Zy8HlS
E0qeq4NtoNN8LwhHwD1pfP+Ezkbt6v7iE4/50lEw4JaEiEHsbSNNEujwC8g+eb1r
FQG9499p+ql1PZG1z6OiXzka7wBGh5JXVHk5qEQeGPUh657HCRzaC6e2TTnGLZcs
dIq/GgJbUCLNQnMJzuakZuqjbMQivDmBtZfvZCrH4fKf+Z04CG8b4Hh81/HLF+Zc
WUxgSVUigQxNF9AJQAnITav7nz8eBiycsm8fTDPlyo3rmYGZU9QywJgd9DLusu37
gz9k+UtQBzffjuMAUAuR7GFFU4MQfpJBtx/ltJ3x2UPeDSuLCXEAhNeEmSzgD82T
e7NnWcuuAKhJPyp615+IMLjWnLqyIsUd/Z232b2JJHsbHeKh+5Do+4wpp4vpRlb9
DmEpaJ1JAB1UZ8gpTZwdp0lLp/GnkqRVEvAlMXkLJURP+BRRbwRR66Ze2Kx/FOsE
GVmw0YEimKckywIblu4DXDyXW7FugJ6fen/ElNK69huEh2d9c5aJ4tKu57Pnp1wA
bt/KDywoLLDMwt35NKu7zACK4tjY0TlsaZmiP2rz1RPgCd5geXNru9K3WFg5ZaXy
Qx9ptro7RDJThADQB9kNAAIuYybGw6FPmlEvRn4YkBJz4KpJWudJS4tr+oLARl+q
dJ0d4rho19afQB7corEZ0+Hf+nepuj4q6bfdj6DUgYaTXUcTT9nvrsjUq+XTqHld
anb6ZbNS3gJCYXAYPlvyTFxVqmxgcYbdpGKf+78CXd/NrtknyVchSkuvomKgMjt4
BNhSYOhiWbJiVcllxcxUvuHspao7KSHxLaHbNXCDxKIpdzsJNOyk2yG0pUFHKq46
q8WQUsbEimXBM1Z36N1ULkzZV39BCdHgyE9ksCrifC7l0hOlWK8yLMCwPa02rhMQ
rMrGCH5UcrBjIqn/ZSZdz3yALMmzNS9o83A2uedvmSHTp0GeaxgxVYmkuUMz20Mm
MMCqEBLjJAgPetM5KbyG7Uq7ZJoEprku4IJgucYBx8pIu4cV6hUCQZEcvdTutcT9
lQs5Hgl++JaPidNbCadUdRWMgcPg5xq8NumeTTS858Omn3FG7CnjNEJe1S64156L
kTfkVscINLEsUuZA509/5uMCil3Jd59ZZ1J95hHbKhwzBDBsvq5ky/EssdJ1uQqy
uexT1OmM0EVYspHafupVxm8pDMCo1xJOIK7MbrOuaCpLI+JosgypHj5/OXvMCdHq
RBsBD2J9BjgRhNRvXVUUAqIWYDYGYs3m2y3BYxwCgVvtkOUOdlJw0O27Jona3jiW
pp4Sdig11x8ZdSNy9abnwXZZ7YeN7OtGk+xHADYzcfs2hV+B+Dz8czmIyT7I/EbR
pmfgThFNy2j9gwndUFW51xUip0j4v57dlgMjYH4zmrTtXgoPnyM/HHe17o9GIWhK
DL5fKuMqQEujo28LGWjRMQRTfj+bF3wun9YpTxnrpYnE4o0Tu8vR4MIlnoaZbpPy
V+jdLwhmu3ltSnZ6Ay/0ezJGfdLeNdhwkOSPIryxYM4F9y3+81n/bmvXHBnwqLek
Q6pITl38nAqM5XQboeB7fHeI5ZE1bkbIR6qN1we+8toiO9Z0/CSekGZD+hWamkiN
EbVVAXYqUYQFNR+nlB+a+bQ8mxcEz3kKG/Kr5TQv4eD+PEzYH1Kw/9RmRYCvV26g
Cp4spPF4uSAS89CFYILj6ux+hYNE+W0U7UqnOJ+1ur6IO1vXu/BYJpjeDXUrXyVH
rgd6I+wEgqvTCRGBNUCms/VOrWIgn6J8N6S19YjAsPQ6S5NwQrDpFG6wI0Vc7NZ1
yPt1EKEjhsMZZVnxANJyjvraP/9/0geqx57XRCCpYMCrAxOOtqHwd/frXagOaX+S
DKeU4S0VZB3Q0f0O4jfPXrQLMCW3mg0OZ1L1PqxslBW7V9yab2lEBqi23v898q+5
apXJScnLWBzwQBDb/dK7FG/LqjF7zcmy5dvupAFVP4kTq4/dJk7F5vhd2SHJGEz1
xH/wojCraWUHcpjcYI4zJqT00uBkSsii+g6PuvaMFE8mP/Y10dDJL2w3YuE5rGap
CFxUsExZALuUAuIYzczD2uIStw1N+wn6YDl2BsWIyxMRCTAcOQ2E29C3v2Ix5gYl
UNWtatuD2hvB9Xy2egtWmjd0N/EErfAVQTusTOs8cHeAupAKv+oDoEKMNZuf6ogu
PH+rwzmEWBZFVRh/tgebGuWd2wDWpoSIbdlmClEBbcIrk03uUoFeRlHzpMnJTrnW
VbQNTC6ZRh5RbYYy0lJhs8StRMcG6UkS2RQ0TsjyNqcb37B3iBGIz6OmOhlS7Ttd
BePvnD+P2A7IhJELGu/NoFMtY5DPBjH4unfAm5572DYhcYFHwqozWUbbuUnwm1Nj
x/d+Nm1YHUJmkNSuW3fiZiP+lAGUF7J6hXP2xNzkI5/vvdNO5tRMkuC5tZmBSSGf
ycYvM6gRnF/ljY35IlLIJAZkjeRCmTHHa/TqPQGuMyUMrTPfbcgBVxwOvkLR7L5j
OB7g9mToRxltfrjcvhD6C2xV0iO0BlcqyvUBUlxlrYeeAe26/yha76OxbkFPdoMN
oBux3h9EG2FAvgFY5Vd6GeqjIdiAS1luY3zCu23iG1qOpBPszBLicCXcgni9IbNN
2I2Skt7lENJ5YUZY9xygTVhhhkzVfhEN19BCSyOBOqBWG6qwjubFZOG/y3PkayND
yrhDCzWHowqZJaOQ9dDOoFM5QG1FvnRLb/u+zvcMs/HIpE8K/PE23aHEusNH8X8N
h4nUsa8YKWnIedpi9MD1416LeHWr9x2TTiTGKFj+uaxtLkPI5g02yPRagkoIxVVm
UBd2dISHc3/Urr/rAbmuwQJmyUgASulZ3m+hwS11rlRFbt1MNhIzHz6dzg8Oimwj
+KaFcPB541ItxkNzE5B1rlBOXuzXOlpAxJIMc4Npc2+B8JFCTpn7IZrMXG1XZsyx
mxj8aObCSM2zpw5GjcC1SzZqo3UF4qaYmPG8TmXjbliMJXnb2JdNi/RafMUOtRQo
BR+auFea3ZbQTBOinYrYy5cPfrYRVAFoH7faqn/ghxujifXTZSGu81H0jNPTz342
Yvh1ENET+h+U6HLQzZP/ShqvF0ygY9OEtdVe+XdjRRqglwnk7GS1tOT1RP6atvC9
X1OOZxSrlu384zZ9kLmm56p+el51itWgW9ThkiFGAqixAVzlb9QG7MrmJ7Niaxff
La9JaURVaD6PK+YcA9RwjbhqRqeTlCpRvcctVC5cp3V/pBDg/9kKWUuVkqMJqemy
jtVsJEiwfTs9Ydey+3dDZzFKBGrMKaH5U194MWdP5EqNDkU89Fhp5O1TPAXn2LD0
Iitsl9J4fWVsGHkp+bqprVzuJwVZNXfBEgFxFDGauJJfy8qWQd9XtMPs3TSPjT0S
JW1wRHK0eibkwWM6S93xnnsym2zk+s1Qrvj1mkOFtehjCDqsAGfRO/7DVtZDnwWg
Y7RYXehn4T7OfxJQaPF0ZIRBEyIIS3NC04OuGxOBCze3DZoTSgXjKeIFur2KmjVS
cD8GlXCpo9Vq/iGXWhx5FpB8PMtYwquHso/S4oAZCgdY/owYc0O8HxXoKpIc5D9j
yVjMFkEuFm+HlRPxqCSMhBdvBAC2W2Oe30fTgVL8XV3nbRp6RYMhGbfNfzwbHbLy
YX7WzlMIHveYv0tsfgmJSHI1oL8x5yeQAXopzAvSqD75Bs5Yl0EaBGBC949ZoHT2
LkPM8dbHhODaiNL5RCP8tG/pm2D7fEcK/CoDom3FH9jqzASIIEuFafULSZ90XxR1
0d2rXW6KFXgSMqkhmLO/7VvJ31rymEJww1HLhAzRfy/OpzvC7B4Y9PyG+x2VF/fz
akUcdIL/lDUrEoOzTrbMngUmHZvNCWegTN1vPFHQuTXEv9HL4QKhPcZgKXlqeB8w
Dmn/eWNP1Go/yriKmTK75r/OMfA6zVLtWpU2LAhty2DXhxC/b+Gtn21ujTA+78BO
NZFEQdM+mzY8Oy9aZ8GdN9Pn3MVEchY+qtakW9o9Hd7/EHIcPPhPunzGLSgNZ5he
H4tJMM723q+zLGU2qB3Vd40WaCPjQ3P+O86MA5EFqBBklUULF5eqeH9twHPdbrX1
RPcOa2LzqE1/qpTL42zvaxqAbIRL9vRRI7Qy5eZSXMKTu1Ri7XpI8ZTzdc9hSbv1
qrkdsyt/nAFNH/G+OXvzJT5gBLif2qgiWWEz75wv4F3rBh5lCrDgfrk7eDkYe+nB
SHALYXIZcxakZF2MWdlC/BO7oJjpcw9L+BB+h8h8cyGhQmnM+y9nvm5yHGp6aL5I
iFp0azFsJP8owLP7vnY4wfQXba37HyG4OPRf6U/OCGNpMziDa363bifuE3TpjH4h
kUTWEmmMT4KeA63hb07mT2j78mf6ecrZMoJ4VxTafQ7uluh9i5BiO1vHoZF7doNx
eCUYdCuylmI2fSGVmCI3xcsIusruzrXL7TAc5LW2SDzrWAdYXgZ567tQXVGNJMH9
vjL73SRZXiusLuawerm5obskCwWLio2lsBsKmv3/+v5Wk7v6eTrzNDcGvwQFH8u3
HEMEida9otDl2cQlc7BJCcHZA5h5qc7oaDgy5A2tAu+mON8g2J12I1P+4pet5JFX
9c3z2EVOp1doMbiTSKsSa7yi+pzqtABKT7J8ff1WKMkn75s0iMnlaFyCp77Sc8Nl
bM8zP9xURp+Uk+0qnvxW1n6w9S0gMJazJie5Ky5eglZRhSy/mOHVOSy2UpZb7r/r
2PY/gtOKZGO61il/mLSp2bNNCgfFULuKuLdwCOrN9n5aRZXakmwD53gIiXMdJ0//
VzN1vuqV8btVnCEAAuOzKQcIOeDul3njVF53CxEg3NoQp3OP3iK959myF/OMIz3X
kZXEPNnnpMpZwqVvkVShf4ULWDTS3t9HqePSIVWCUF0NA1RhmQ3S1O7/hHF/Sc17
MBVb724PiNc2lVoEcAxIQSluHGC29cVPEDA2YlbMgl7AFyvU/shO895pjpn/18gX
QO6FNVfr3ohyKsWKzTt2HklOcpArlejnTXanINtKu+zwlzKTysRU22U4Dz+GxIGZ
VYjCltf3mcduMkCNHQfFyX4/UJAOmDTV+UbvIGTK1gpZqHFdpFOt79ythjrXJkUk
Z31su8X53TouhkQjSmhuVooKCyF0D9ix4ITSkl5ju7b/hs9yEu7t1KQMlPYsWsbm
lq7dmsR0It70AIjw+2bscFHRtTgBmghsgDvhBq1A2DLZrvuZwOh+OeqT+aNzMDQu
RlZIAc7f3Afl71yE6HYmy94mgbl0z6RdCxXfiMTTjqS13batS3g3PX8VzjJVQIZN
z4u4GExsRhq9Ud/9xVjCWrVqH3xRfOsEpyZUcD7HtdyzxlaCUy6YEn3brtrCcOi6
3agBB7hNHdG1J5LqD2cN1m05nce1BY38AN9AM966bQCLx52XLhtqP+Aeue6RcVvw
D/BQbQhtr9y0B/KppiEcoPs1B4YEIO3E2W7GeN6rF4vpszw9ZWl1eNKKbZt3z8/4
CEVce2aj1tyP7Xk371NW5CWfwjzGx3mUx/1NU8b1CclEOPG33ywwY4NdbRuhWi69
TwZl8pZS0FTwQ5j+2CQGnLka029RVPMl5G6n8FQE+3acsBhZM8C77E9oH+WU8IzW
ECIMg0+M1wUlp663pterGvBGQctcAdf3gDcAk1MIjVmIQbB3+DiNGIZtJUlVfDPm
bBHtsbeSujWDnRYc9zJvuMwWiPcOpMFXm0BE+V8jAdwbyKbdIrF3oNsgyoFAohtg
b2If9xFFz7dYI77U5IXPrGpV0Xik42lTWGWGECbG6fXm/Mtfgx8fPzeNgB0xeLk3
pYl4QFVd5U6f+RiEgkbyzUpViQVo0xe0Ws7wbbi1tYbZigd9iLGc4VHo8YxocTFU
ZFhEWV9VbfUw3t4M05p+6kCZESX2sUoQZsLls4Xw3zESG9F03uvK8YNYMsN7hp1X
1zA//+wY3KfgQ0kGQ/JWnUkzmOFuKJUif5iw1xlUJa6FtmJe5Yq5APoI0o0tFwF8
CziXTgET3Prf0FLOmfolhY/GIF+GQK2s8D2sqWdBttGIZBwBv3ft8CyIwgIVf+sc
Emb7CK+4teSNl2Rwdac5Bjg6wI99Ttya7mi5yuyxjRPQdseV8nSBPiXTKPAIHGI3
MqQ+zk09LsTpcAubXtWqaMZN9sL7On6TKt7lHpu5ttRPeSSFqsayo6QbXWeeLyxA
m25QZBG2P9rCtq7TV00RWW5UI6fD9Er9ipVA/1YSPnoKvo1NY/3MDRlWG4Hcb5T+
v2OdVdFZYRVo8pHGTRw++VhwdrYtsKx0EsDmnH7HQRCktX1LDNoonnKC9ObhwC+S
E3JcwHCsCMDZLhJQRysjNrpnvHgEFrC2qQ2M+AdFhz84DZPSJ0bXlalRm5kCTyV5
Uab6mvOdGdIZI++pSMS+VO+nS+DIDrpBjMosnoX2L3hdmw5gJqgTXe6Vq1qfXMdR
DUcYiukm7w3nXij6mkFhjVgTP4xnM2pGqh0ob96yH1PQTx53XM8nKW8dwZYNTPid
JysQP18P526hVYHnFiTao5TZpE/L2tJZ2gFUD+hcRKpSG8gM0AsvraIukXsOJtVL
f8arrL1bcF1xRJP1UkRp+VnlAgrRaNhXXk3fwg2LP50UFG8y0g205PzE2bYcj6LA
L7BMrZ3sroxmSi2OJz/9o4vdUC0EcM9/kbdBQ4c2cxUI3fB5gYVcQx5XVObpBkhl
Kt+jewmnQKQQKQI1AnVstUjY+utRSuhe37aLCmUSZIt873S13cJGTb54mQ9uS7ym
T/1S+7o+A5k5NiN37qsYOQK8miltU2UYWezJlW3DQPYukOFRvqzSL5q738mfff4s
XenKOiYB+uQHvlAdme/DxFOdLxMj+PIukWhCgkXJPVxsG5UnAb1mY/TR3aRuN9ON
uwAgQWAFerwAyyTWD+iHf4/34S7AUWSD0YUrAStEm6KrkH6bts6J+pz8uZi8qU/a
zReeuapdYO2DB36wASycg1fOhwG9EeInddJHKFnAaJqNLn1nTiMT3PpMPloCnR2g
1AfKQk2LzEpwt7RUdAZpesYusa3f6ziOmig0lrGwJkCBhC/g/fPGlLkC/G3yKz+/
466thjHW5Qfari4AmgqEKMqYGeL6JZltSo+/cjypPKlkjvvz6NaBtcxxA8X/b5WQ
NrGnz7P61j6ZcpeAM42hcSsaTD1dZ3PosXp6AFsMBpPn7due80MGAZP/zd/nK4eF
5MJjvdMnBJ31ljnL883UCvJrQXmR5lIHqWfb8T6EkcW6qwQ8TJozYFywQCn/FYaO
I2PrEp2FmSO33NQHqH3T7Jl4iGgxhfpUn8mX15eDw7CX71iQZIPikOy1nD62ODHH
A1EkKVSPzuR5tIU90I0Ed42qihHnKInl+5/GGRi1S36knRD6rNHy+D4QY8+M3EB9
DFeQYXaa/jKyFiLugnKzgEKo14EGar64Mqr4WZUOotX8k+Q9BLIYkaOgHAf2q/Z0
kVAINZAk0H7YKpoBNBbCvHwbfNYrqo68jBaWSxY5GFCd5k9bAItnllBgpvkKvy43
Kxuv9q2SIW+kjSY5DeY56zggC0Ful1M6W5hfb17P0sQz/uPxCs/20m9/hbqgW8RL
3PWDHsiYWpkug21bEZ7oPqph+s4tdFRG2cddb5SwUS0ovL3EMAZ4LRJNchvTV3BS
FmtJjViTina4rW+Ij88h2SM/9gQ07XicZ5n1ZYQ8iDqJ7jb1URV6+KttZt4WWk3Q
vfx+WUET55rzrjTf8e7t+ilALRAV49MDOWTxwWcdguy6GMbP4SyhjTc77BrpfxuF
X9Pax/T/1++DI6K9j+8YKJgjPUfAYiUGLECwFSOlg5haDBtKgXAsoC1iyVmT9H30
wSZLTOZ8omi+QS4/pZmkNAHSedu1o9/NrFJdhbgOspb8IXDnuCoc1nabWBOZSlfp
SmLW39SrH+p55nwYcZWqkhvXPA2Kw8rw8G3B9rxLusFcm4YvwrqKmv3d2wN+QfUE
NaIGdUHEb4gUEQFDa/34tsNfEgwl0jaMZTv4f4ULprkGW46tLo/icbxYz7vvYTp5
76eu0HJ77FG+stCjdGs6qWG2ejXGHd2zyhM8lbQO1wI1yRQ6D3bsbGaecL0oePXH
/Ni/h51JK2hGinf6jkDqSKSfunVheIvNEAcMWOOhjrjmW51wLw3OhED1UwaF3320
ceZyjWwBAe/bcOAUZIDWy8DrhaxyZidwyJJpM6sB4j2PKuNNVeYtcQz5gog9Q1Xg
y9f4Vkegki3dDdsN93YBvThM5cJ2ZBRH7uTJmPMittkmou2MLWvJUeHoR9SMe7lT
810lvIpU3AZ7Hdrr53GDC3ZM/JwUrrXrQI8Rz4XtxHp+3aYGzO5lRBYzAE8J1fqM
+1AXVj+/KAL/R2r8aGKcwfalNB7B2VE1xPyfM/luOuhil9mslg7lQg9rZ3LoAwPa
N02TyazwQTGBmm23y8NMZHnCxEDeFkd7lFVhEd6Omku8NORaEwQfxf2Bz0Z0Z/j5
XnJ13BmYzywW5sPe5HlG4eIiMFZ79eGU0sETKdcLTj86gnOaKjzYGF/4BkfNyzjs
03QsXp/aA3HvpAYeRCMKBIwMKA+RdputEHNMM0iETRgOuxXGkBembNT5Jpja9dfN
PSoqvcI5VP+yQgSPYcG4XsPzCmk3P0X8FJvIBDt0CUM6p+qxJ5DX8cCecwzFcGFl
aEVd2Ib61jXWHUE7vONxQX3/yLQp56rlf3Fw5787yeda7PwNHcQcdI0VZ21+MfTC
MMUUVXTjLuk7NisqJ8eXnGfrssTx/DctKclP2mcT2fRV+ukBw164/GsJ1dVTsbf+
UipkuTtrKHq83F7OM51okcdUyobW2727TABvuFDRUEf6alfUKvBPlumTH/EpjFTL
Uc4AXwGRqdVil45J7hZIkyLnCjaxdWS8YqVrwCj/Jk1O5zxj1B/CmRcLMvZHgGbn
Kt5RtYY+4fQN6x+Q9hT+9H7FIGS+4ENIT2KGZPCJK1wVsA5QfSY3Y0UYOvpOURqh
kSpjbVBffiyycHVV/ZXYD7XLwoPFa1KP1N1b1klTcycxVt9J5Ioo90xMW5TCY4Gq
bNow2i3t+/tDqTil5TRPwauKKg7tjjGiGiYPy/TftbDs4yaIgEozvwvvC3nvqn05
FHT9FFfXFdNmYby9ONv+mwpCiyu9kp03rJ/LDbWyj8/40RoKksDzLCISVvDWuath
gXtZsBXrV70sLZSoRnmw/j/THKgPJsfOI2r8ymKI1wWI2hzCvjkSaYKXFsHaAWov
XqlQmhywzbie23q7E+e3Xd59U3osLbDqlL8jFcFWIBcqWdMY5BEHfIzmvjwDREze
r5HjYkvxi/Sp3U5WT9tj45MWpQcg+7GCDY2IHQl1moihGf9kTkZYGBDmkUZoHuv4
uR+5VTIfNP48RW/EMf7omrd70Dxp2WHy0E/LsAJqCzwwhP1D2jAK4bE/9/TC2LD7
exWVz6cg1kxHhcY5rGtEAu40apkplAhqraI0ExBgpGNe/rx9DlWB5XG+k0K7QrRV
AzEhzJED+BTDvoDnZmWTGDEByInOSlTKL/XgmdiUaXafgplzI3+MA1jI0lqgufws
ei8h1+RRXbnGElBU9OQnWue7sE1/LsYpSWmphp7XnuGcXQiLnunXN0S/uPquwS0F
AZH2rIRfPfxvWqfmtNSr/KF2AykFHpjrdMVEZKJm2pMnXhuoQ5yjNRILwEjfvAtT
OVLuC5md/ePiqdBYrFL+6CUpxhOCr4lboNftmzUBh2B0/8Xn6YFRQIWhVjUZv+6G
lr3ZNKjbmz+ISn7xxKhNH1dwbo6W47kWSQLBetPcMapv2mej1agDezknhw8aJZ4+
2w/diCqBYVLNyklTN25sM8of2eVHjcxFq5UaarsZ+cDCC8aZZ0Omcvb9kAPgMXQs
8l9NeaLXfg55G+Kksr91SA2eFW9vY/ifeqkUwL6ucR9mTTEqzrtK5C5PbpjFJ5Z9
SkYgv5SHOg+HJUL6HY7f9k45n1BKzZGq8tszisourdlhAhbU1Dj70jePw+Xn3iR5
OJaoosKiAKZXxs4O33Wom6LbRFNXUuW2K+bRwFtkVPGkyfLA5rFQS0hByFSnn9Zr
C52hnHWKhRJ53KGgUDjD9FkXTL/vp1/dLxnXNzrRkVFGF4Li0wnn2q1iUe6T6sGZ
Sy/jjFVWR4nYjVlZAmAh5vkZs2Th0+zKRl7TlioKXwbsYr+UMdVZB9CPlafpSM0Q
rR+s6aZYSZ58vYSyscTu8f//12wIBMXoGEGVnBEHKSJtusHGqcYIYJVdj4OVDk1j
86E3SwYqaEQOmZpENcWJXhG8LSYx5XWIaoXZC2/rtiX3MGZuWLRQooRnXVOO3QqI
6GNXLXxJt+sKD0uBpZKSqN77lsmUNg6EecGoeutj5hAq4EvmFKiHPginG8SFnxXy
6r7CcYr147EnAcZjmmCbEibkd13Vs4ycDaKNJ8qUWrupkROTC3bDJxyO/7Qp2KAn
BPgQzniFkNLl0RH+GdRnrRX2g5yLNa5SGRycE5iDWU8CszqEteOu6lD/2IvcHaIP
M6CH67/irfpz0Fr+qX5gA6WvO4UqlCp9UAarPsRvIKtTQ0QzvAS5HXgVnqb1AAEP
kLjO0fe3UccUNokcE5LBZLZBuy1/ApS7F2RC9fhoZjb6R84+3xsXJxBIlb+ZAgV2
bNCQhMOXw4tKYwyY8nQua2CBMGQ08JXFkK00HufnloGQTYdCHMb467UFPfRYf/Fk
YsGaXO50fdESJVng7FbcoygXZiWzyvAxvpIwgUNIiBSX1PS7m94PExnjAG7duCqr
6ziooz9OGOTx/1xi0CphCJDrE9tMrtPZkb71pFT2XTVATv+YYqBfzvvjz+G0Ntor
qDXiheRYBA+qGT/IdyTGKLv+1J40cxpmywQDHBcbE1pb1eEFX1ie9E507/I2/bph
1WWV7qGiFbpHUEh9EmFz0Q7Izr3fSpPruUiWrmv181UnD0p0VuxYNCO+7wnvhCru
b7J3BcoCvwYp0L4BRxjU+niq/QazZgb0rvEW8QgkKfRMNda2URhQs0zL9wgYHBY3
omrzEdzyAFSQWZICgcg6+C6+AukS9j9hjHlwlIeKlYCkR6HgR3T/GJoPz/005WFA
mU9fUauJ29NqDdblHlk04g8iczjj6ztsjP3QLN3i1nflPupVr4hL9FHa1xf8bcPU
xC9cn+HmuRCZ4mKv2qnl9Xyk4vZWhZxxb4BYi4XAUC52AAzZic2HJDSQk+Udz4eZ
xlyFMM7MunJPSdkIeyVIH/ywQwA+9kh0QLB0/qAGfJjrA7NfLR8NgfmuyG2ul9/3
E9N6i5s4syD34inrYekQL5r6HDK+IXX9aTzRh/A9eQmdbNKQq04gbTe3iScMZGxs
rWRXHysCrvH5Nk6GOhsWEYAMu5uJd2unKcSmbCZkqwBfdvK0bW0PkUATTGVo0F93
hLgM+SEuvTUVqToaEebOJ8wStJNRSPma+KApyjgpQ2T6QOrfhcNrgE2Psftju8hX
mi5l0B/9LMwi1IGxJwVT2cNXIcyp0nxRc2aNCFa2w9YVtvoh5GggXJ9PfezHf41+
2MfUxB0BPTkRsNgBh3oxw2I4vyUIiJAB9d61oZ5Gw6yVUQPdupQKt7WZ+WkkcLbf
5VsryqFSqUvbL9cAIT8bBRzvXJs1M9UfO8ug3PN92a4IBYJ1UB+cQ4+N4R4cb1/S
awSnOdh4NB5IBk0B6iZ9qSQ9MpwWcdzVoy31fDlH/9DT1l4q5VlQPORLmN0ZeOIf
KP+eG/HAxPffogsK+AiRXogU6ivD0xPYrjbY2HdwxrYNlf3PQfXjaEgq5lOKbLax
AUNKeHnUH8sGFKqedpwttIrXdjVAJfeo4JnW+Z0NtkvxuJKRz+nWJ8EMxcDnO396
HhEUe+0/P19zSYU/VI36oSwowMxdeMw8VCgTXjlfL+FzMQ8p2zZ796x1CIDFCwil
Yn3BLdDQ6ew3sthA7YEHaW0GvYBBwykaagd7scU7lfycL7OW64/y6t01fzO2XO/P
hJdX9LZJaJSCK20MM2zmKPAT4MTqxctJDeiCw0VthZ6OG/J+iUje9v+UYmij+63y
0veLifiPdZBMROAmUleKzLUcWYVhV7BcwDuzSHDnYHd+4bjMUrobYh/j/BXd9DRg
CoJNtI5ZYFSpipVdJ7r8dAfm1d9OOXmNliE37V2dp6nefiihg0rP6RNLmUwy+ukP
RXH0zNgPAyymXKhlwfadHgL407YqzvBvOAinfFynxWbJhyZwUINLWuDDw7ShxgI2
jTSMhaqbA89DsZOnl+p4KiQo7QY4XGjjzLvwQRtE/d4wjSi+obRLP7YAwfeEJWZg
LSHmG+syYMdhaHcYiFzkSiGP1OsA1URLW47/WexgyvjmXSmGSarD0dcElLSHWFlA
Lt3dHR4RZy9gat8Sa1HjJUWoY4u+3kOiWUyOzYbHZz3+wtuvKk9zfePQIOPcVIko
zq0ygBsY1CmG4haWdgQzOMv0Om92S8lrSi8RDs1LUdtoe/Lkxl/6IA+yN+Xanfpr
yWbJkyQFhQ1ZhD0c3do5hTG5Nk2UkIPDVj+3pBoGCMOMtRtLPK6DtPk/D0o8WsPp
bupKJpjNb1ALEQQMXah+ymR794rMXC7aXDtLAnKgJCIR6ADnMYBcyB9KMuKkqMlo
5T3R5ZDUKuSlSZnkBettBsclMxjsjtLMPtay4zgHCWVKDWy2u0j2fs+h31BWKBTg
TZik75q0MPLBBFo2lZ4MxLkxWvTBRCNVNlnp2fe7CGiPflD/PVQ+7uUphXKOAy0V
rHQcss+UX8Vj59Ut7m25g2vV6vV3cMO8LCw5SLnNiVtfOsaiQOeCuKPzxbxntpuw
VubXfOv8Y+qtAfLywwPpXBcCQ3NRP7LhDazL6PcBuU3lMJzNSyMrZfhvF23dINbN
EXJg3zyqkC3g6Myha8N1f2Df9vTi/ezoQESkrb3ptHbTxgCjrtKPpLvpG45UtGiw
bLfeEyIzPTU9QgkXszsdbykutNYp/AhXSGe9bdSkXoqdh9rs01ADyFXa/mINKvR1
qzyM6LXf0CWHRTJ8DJTe09qTn+K4iyP+M8yRWgo1y0RsUZaL9KL+IVMhtt424AuH
3LtmMO7Ngcx9bpp4o4Ae/VJga3Afr6G2M21YI1zXjrDSfviqBycpQxgvFfPGddqv
GCpHONWYxvmbA+mYHc9FguOc8vxM8Dv8ToH703wibJqb9dbLUqXuVaQg8yOZPvi4
keel3+LLVB2OxNM6Fbw5TG7ppdkIw+rNmYOCFqrrCpw8HGWReAHLdnxlXt5hUvET
vfVF1n1EUcsPE1FkafdAYTcJhwRaQFXDW9ut9/y7j0SquD5i8reaN1L8ayZzsX8f
ABKyfqCmyEQNlHEa2zGnuhZdqa5sy4vmIiR55DUO2+zoVNTAFuX/vuHo43Ts24sh
3iD9zBRnW0RzACSLE5n7sFh0Z1E2Gd/QNBwvgI/dssL7mp93VPzWD2iGg5UbtpyS
D/ExdcxxHd4QeuA9rCCXjVSvfCVIJQ1mR11Rc+Uj8zwVq/rYDwyC1cEdTdBtF5kW
kuRCPlHOLDGYm9f7biovkoVaMgtbVGwF1IrQPfvUW0bPy8dGARFB35WyqQEvsoYe
EPKvycjMl4jO6bQyn4GZ7USR08Bk+ZewfF2NR0eKL1vbT0IIJ7ERvqa1D8J2X3ut
JKo0zq/rE7oArriTAvhAroFd86nvHdqBQGE50/T2ANlUtIbg/hiJjIqviO/GUqQT
e6HX5hEguhpAQ9XCQFU+7KgYTIFS1A2FAN7AmIxSnQAIQsG0+Ot4EqCUzbT/07JO
sP2zw9Ms/31vwpFfRhpVah+yBDnnxo20CHNVPqcDDbQxJUxBVMydiHpQrDNe786a
KWGEa/4bJGN4+C5ssrt94FWkPKV4Mccm10qJuP3S4vYhBf9+XdgEXl0mA4PSfrxZ
kkrTqg4rOmYdUArP81bBgFoQDs7KEHVKS5sERFvDjNFHCq1kJf3M4vBnkprb0ZKR
44YR3CXHNnHVg8LvC6z5hRPmpW1K4At3FJrxNtmJ+tvw7G9jzdBU2PWXarzLz1+R
Px/EUb4DNvZbDFLR6sHiOZKd+3Hhy2g4RExswAjGXnNtkKBsK/QPusnXlN1N6RBG
vAeQdxsJEW7ZYI9t8eP6eYRBYdGDxUVUQuBeamiYv2bH4CVEwuab/9ai7D2R+uDA
5pwK0vErRRbSO4VggXPtaUiwMG20cDPSCJlQlzlRGwQtcHTm1iyA3QjtRR9LhgKg
g47RoK4XsgW+O3bEh4YOcMIP7p+EyDyP1JYOqwrxAa7GflJUCwIdIg4tqfHK/Ubb
ZhOPSu/h91An/e80lYIomlFrTw0FLn96l/mg6stPPIGO8CV+A65T+U3vKFp1KW4V
gkZ7qNZlkgNvPru4zHOb392Vca5FqH4mx8On7ZokmSJFtA7eGAPi7ofXW0NfXnpE
G/ZsPMDuSYVqdfkx0OGHuwjbHg3R2YRAXzo2aaygTBQUVFQdVf+KlZynzEBjUk8D
8Bk1OqIYd6nKWIHvnR8UAjBqpC1yBWpIfJ4cf5ZdBNHlRqmH0sx3hbHLtDqGMWy5
qrBcIX+w6KMoISwKqpN1f0sVHe1G12UCLsjLybJKu9thuX2yWkrqtClTgEeZ1+7O
qFkiih8nQqh+/bDRPDmQC7Y81e/g9P8ErgT+3a5oHjAaaSi9Qfj39msPzYrkECfG
n0/jjDXFHlmB1J8kEO60YX2ZNjoox1/Cqm5V1hSThb4Mp4g79hrP/kls2gMHOWcz
KwRU1VnYnyt9eoAb4jtJwSBVB+6CNlWFXl5EnLfdRm4oZDt5uAXgslSmY8B/yXyg
MgBT3kejdVoCH4iAmD51uCq381Y7spLyLGPIOBw8fy2Esd7hWb7YXjyga4SVBd13
af3gTSWhGVf4OGFoc7yNkjXTQG9tarh4K3bYfHZFeJOVbq+qfNhXKhNnGxlBfHGn
sN/hFCN7hZKxOfXW6db5XPNCAHCj03nAs4eylAGsypcDUCYyPNyAZDGjbnXcA5CL
YklTy/Jdf+2oetS1Ax6AXqlYM+rz/OWrYr/xL4zPVqdMWtsFI6Mlot3jRcgmfIy3
awCmRA+u6NulSOMeCo4FIkdugubZBuFxBxZDN+lHyS+Wkyi9Yo8YGq5lGYUH/1dP
BoWK8s6SivzV+qdScgb4XlvfdbS9SFUophsrDTxwYp1sFo+6kpx+gOvZn3M0NN/h
MRNknOgo0W5SNNSeerzlWiAJz24ybcN4bkrqQO/g+HCpf2+rbjKk5mCL+Xbzjo/k
0Rkkfdg4x/0hvXBTijy+9jzIU6FrRAqL30lxxJw5fALgFbCiBKKyAf70q0Vo9rnq
ysg68Tvt//DrE+hyl6U/vc/V2lcDZgBpuTN/dStYNfdv81Kt6oU/FzZdZPv60VjV
T4DgdinVXeFHItQLiIobT2J8e99b4FF7zdIp66pHOSbkP3+qQdlj2ro2CAXybKvX
9X0d9KKEaJMVi7OJOk6/Rpkq4NIWcFDzvy2t1hdeit0psJbmvNrbU8RxJsZPsis7
1AIp6LEWX+2aqrq7RCUErSJoHDU9X38OmodVNOVGs1NZqNTKsm2w8GLJl7cGKXbA
uD4gddWeP0GjlTRtGUNTosH6qI0nKDovt9vqgDGoCmgFNTPNnw197f5SfII9TSx9
qPeqBrykyZL/8gBOYFCM9Bsrm5fqKgAwfcoOwAONWkQ/ETD1mVVLk6ptcit0zIpw
XHVL8ON4Qe7V6+K3jA+nzcWT3Bdy8naEBPN/if2eXhM1inuLtvhEBEKgrcn+Xt8/
ku3N+DsftAcwlGIkZBul5rTt4xoYlPGkgJjj1m+B6vnjyJ4xDU2fl2i86/pFkMf5
QjnDukXcV6aGVLKUq7Sx4MhReXzlu766YW37fhgKaYJgjDgUApdkI2dLGZE9DVyN
MNviZXUXCyQFu2RcwkRd5qKoNajncUijwFiw5XKWShffs2lDTGvOgkIRexxW023M
p4gQZGVIuEH5I5ogpvYPmBNGoGCC9fmIxwsfm418TMPBwlMOkI3xorOghcSV/LPu
PrSz+mqXVyZNOzb9OhEpu0ohlfDdGhhTuI1jtP0zpUPMPPr7sXGL0Sk4VT/8eCVp
LnnE3Tn98Y8zuZJ4jXaO4lX5xxI5nItEyyp74H5qJLvrXcL8UgRyd6yAYXbnIkSb
WI7OUaBpXNKrVVqelmy2qf2gCas+0q5q7CZfrPJHy7vTskbMw4SFtpW5qvTnGJRd
2YQvBxQS899lA+kopRjzKE1auzHd2ddOwnI72Vo5as3n59/LMRt9dztF8nnIFUeb
5gREamUfbp1p6HLdpahol2AFn14qSKNET16YU5wgS0ggmpZGdDEml0LtVGbYHB7X
VDoy3ewHFU5GZZsmkb2ksm928jN0B+lhHRIT8cX/aN3wt7ggLI5nyPRrvWX5uFd0
Sh3TNNUEDeJpj28THf1WSI+Q2agBBG7TL7MHJ8NBsGLtM7pEMUUtjKl04xV/c2mm
IUCUdFbZq33luwcnpeEN86QoCr8Sd8A2RgBHuRH7zRzE9eoM7jUdiYYiHAmspU/T
J5ft12/JcUWtzzJR5tUEiCpUgnsG5orZlAbICkymp11kee5utfjHTlssD1LGZwo/
AnQwbJGnCR0LTcxB4jHFSOWtAhRgdzUz27hZC+8nhIl4d5bqL3Rn6iKirNGKV0NU
L8M8437118Ow6xMgaG5SPvs8mBxlSA9HOboZQGQW1MDTnkoNHTZejy5/ntxMmddg
J7+p7LqVKc1HaQlKqD3/48hORmRp+O99ZgiSHV/rcVF8tPqr994tXrKBi51N3U86
YKNQzVb6BfDIyfy+zvk1EbbQtP4kNlZoLgyfz/VKsQNC3gAMJVAMmCNHQ+aZ5w6L
LPVEM+csZ5RsHnXJs0U3jO+hJUawsVRP9QoqLt+l4J9wZHrt2z5QW6rhotEsWO4E
tzICN7dxzKOwRXS14gRrKnLTGV+zQkH6LnRtRTXLm/vCiI5pGTLRv6UnC0RavnDk
Ehm9OMJm7i8AETNBVuvXXhVKEypuEPDiSX0AZ1St9K+txfpv65RKMBLjkjZ2SEQ+
xfkVxDvPAkN16pWU8srwK015lalFWp91bd83Zhv9pJm9zWJr84bRCPVlJNZhGWCn
MNBvwTVP8Qn0X4TEMdeQl6O8m8DQDjhfx7o4tPOHvB1Y6nxHoXZdEo6FmZ/NMQYE
ncOtNU5geDrpbXGjAtaHccP6p88/x8XoJc28TWVmK50atMbj4Y7rN7G8ufTJu9B7
j5R1JyKXKuaFaKQEu7A2EVVNtINVkk4YCUDWqnNYX58OH6eLVOC2IDCYlEXI3s6R
JrjTiFGZyepBzhuKXAUE6eS3XW8G9x1BMvpcijmR2pehvZVMxrjSCIKpdGwpcLuo
oYY3URASPzpl99UaIr5GE/FZEoahkOpyo/rrREBmRVXFeOC8efZbkU7gRi+WOZ5O
/UhQdFUnTgUb9kwL8bCel3io3WPYSAYC+RVvOn9gyJzQ43oAuUqUkAan62UYPinm
+AJbv9LL1Hoh9ijpgpNarygNlH8730nSMEqNL3KMI6ByowMGHv8qv34Wr8sw3UTM
hX7afKWl1TawNMdcwB1hfNC2MymytoClfmH8EkPebtaSwKbAT30s0Q8yY1miLmOb
lI1A0Plt1pBtUjuloO0qqf26kF/Pud2INLk+ArclMsv7Bnjo1MjKE9YMT2m9FHlN
PkghSeyOcaqV2Wrp8ITouClhWm7HnWpT3TTFHiK3pna8v68CspE0QXo40Wt36ZD4
EVIX2JZ8brfBYGgL2FCQS2rvZ2Yh0DpV90jMIKKNeOp/DlK8xKKT5IZEXywVR/9n
nSJXEuxLiE+SbjKVoBl+mph3J/X8phxEixz5u4dY3mUi3GrmFASwcahDcQD1AZPW
EcCTyapHyvvDELpZKhkOpCBRnff0PG1koiAPqGb0NIp+P5SRvbTjxT9qyZG9qhmX
dxJEaEbaz4SYSZMcVoTOz7pZwkLG2T5IECHirBpjj5k968aO7LFSO1K5FZJrLjVm
BV4tTQ1BdX7O5QlcoB3e5MMdbckNsgzchw6ThjxgoHWGDhHPep4TrEhElHQll0BM
+TX/90rzr0vPklOqpLwFMHTHN9WieA0vQGOacBaZRl2WNYu1pa0C+Kze5GaKLFjW
Z533+jRuIyl9n0LvJNULRpqcTO/McgYl7J/AmQZRnbPAadfoFmWK4zEt96WlZr+i
TfWRYNkzNf4jtogrFwkzXpP+Y512mrX32J57VIffkdn0C/puJ4FH1bD/ectdeI7z
vl5hERfjVVy7JUexyIuRLhQxSJCUPqYqb3j98eZ2SdbuCeTrXyKIuStzlWbS0jYp
zRpsN7eWMNiareoKrO6o2GOzJfLb9D+S7bWABdxN1hI/y/bLAzXQOkuwE+F3qVls
JzbDNx1mH0PQ/4kp9ryEl4U51eXJPb7ij79E92VA73aek6YDlv2RlGT+DNztdYwg
4gwO9vIqUsOTW/b2G9UN8YyXdygao1f1J5t4rhTUZ2kgcOlO4oRHRkLU6unkXBCf
w2byg4VxAyoGj97/Y0KwMgNZ/solvWVIddPldJy2dGHgVNJVHPhBu70YsDTOLafX
5kHghYbV1mBBANNKRphjiQOztrC7za8DA+FUkCEyD05UUNvyfqbKumIsUc6hBBvc
nyT1N2W4uXUHarFvW8bJ5hKriJ4sUvMBGYYXByUWwxlZEe0TsfEGQ0YluAn1TzwY
TBJ3FouASk7zC7iRLf1TF4Gtg75NpwU4i6tHC4KLAuedf3BcXek6XqlPHf+p6HwW
bamM24r6QvJxp0fSO2QO+uN1tUinQsVWPGyMIfLqLx7ng5N3k4abcYGxp/dnpDFG
J7/Fhj6A5GvB7qZCAdNseSwBLQRK/4Hbbs8ZlCqghIpoZCUGefed3RONHaQgt7Gp
zJ10dddHF6nrqfjB2dDFd0moXdfGTJOL/3NrE8bHSxFvhVxLYMwfAkwmTrtqudTV
goE1BYU1TNL9dbNd/NgV9VFenAnT8PLej1CitwVOGMxwSSqMXdxy8xAiF2n5uEC/
2J9PyDQB0BqjLMvPnqZjOEPq4ODeUnnDE//+mOpo3sFRajYqB136fQmYiLTNTytj
lS9oIxtiiG45LHi7rxN0OF7AmCzUD7SmlNvbHCq3/oX32MWlDUq9+/BuqdRg86+w
0+7G0XDdocWbjYwHYuQgt4wk9n4wjpQiio6LcRiwvx9KAevKBb+kmJWetifR6HuR
U/wi/HgeC7JFTghddjmHpS95gdQzokUacE4Ed0gL2xFnVDw5P/egW8E5VnK08Gol
Ul1bcyElYh90keJKrouxyNeoxENcgmpm7b/G3CJQ4u2537XTJbCE9Tx+Bm4ZL2Mt
/elDtuI4pCN9/U4oUO4XMZVA2RYRDgoRB/RaipzmfZdJtVkoQlUaPl0Fpk5XnLGv
BGcoSaJG2GXcarACm9UWANFCdF84wCpIqCfZzhCMLPxK5+axHqhBt/63RO69+tt2
YBnmJ4u7lCdREHxoaI3U9Y/zpzOheebPaREp8CfITYuBR14fjW0u0EBYYQGk3nuR
cwZrm+Qwxn+en2k3Jdj6LsEToMmPDFmqz8FYG9Acvl3x7Je5TI3OxPmGVzkpqksf
kg6KO2e4dDe5zeM9oPCXsM7B0CAoIh/me2rlLx95l6jpBi8K/ihTtoYA+VgB0Ulq
vaiE5j2546HzOMChd9pWWzYFSTN+3SME6faGwV4H4qYtzhUvxmi3UqP3mrj3yiOS
Y64xWHAF/cGIECoB6fTWw4mowd1scNX4g+mrkb4Rn3wZxwJc+zFcU/TcFY7GS6rt
kZyR3x4+Dr/smBhn+PJ9UTub3G0Lwl+wKzgkDhhmh5myQ1uZyWLHjs57t0QgUzhh
2WmHTx8uQNdEPlFlpnImy8IyGyVzjSFwum8INUDxm4D9R+b/JuDC9qEzr4Wfp5Bq
PqBhR8F1bHZ5DjQVX0N9YL4ZszHQ1/Gs8TtgNHCz9Lx4wcLBMQLJytv8ze7Y7A+5
u+tpWYAIiS+tMiqOcvvQuzbmbASIJ/bMQSL9ZN5xx6/hR3W4UrnfiuVbP85JXJrm
JWyYo6AGJkAXwiCPtTzlZn67I51tDHDHUNgeXtXo5BBxljW51xdFY/A9MDb+YN/H
B46pjYkvkwfyPki5M4JUV28Vg9sfWRRwop1Nqf9JlQO89fXaa+oR4C/KeQe8obka
pWLAt2GTwwM+C3zVyc56AsL0jZYEezJN92IMrzauidbERFU79Q+06h1d2Ez/qC5O
J8sij7D2uSYzMk/9lR8i5kU5UhR7nw/uz0P/CpKurF4nKQAQkOMq2UNp+hwfPGlm
TR10a/V4trspjGPLCexG7q548EGzb2cxx3b9TfQhkyhojT18dh2JDg/HLRbApaKq
UTHqBo0xBdpIgv4YfyWr/CtoyauTr8Ll/U9v1B1IljEW/96Ziw4NMdJcB8rceCB8
RUola4iGnzlxUKLbl7OBLFpWR+Q8MPFx2hlo0gSXal8IA8FGTByqNHYqaHfb/hip
spUyJEvtfvw5MsiHGgTdtXaElZRWSUleLV0Cu9fthkUPeLHkNygAdmQo2qU5kXKk
ruoCznYZhvDzwjyYa8sSE76J8ntDirh9Qt0zr2ZGbgw9bd/QGBGx8w+8O9vxBNNH
7e8MQ1NiTXZojjxR5qyVoSabylJixezrgWFaW4FhKQhGthgLxlPNIm4IAfUU2gRN
hvAZBIwxg4ns2eBm7P3rQSNMTCN4yJYe5ZjZRsJ/g1bUlO4E3JvIP1/TRpJ0fdxc
0oI0G9qqm3vxrkSXKxpIDV0z2Zt07S8sZA8uIRBUjbdYKAn4V48CXfqA6PoZbHMq
Azw29CAG7+EB8c44r2b8DA175jVHUlqh8t4wjrkJG3hHG27vEMB7PIKfq88HPNxY
rr/o4kD0pKRPG3/oLW+kRUqHERS5jxEWehnj1S94HsgV+b6JR/+wN89+eS7jQoBl
/WErSoVL6PBSroJ8qhqkCXTTQykCY74xGaKm3bnOBCKgFfDdLba9zwymf4VAnymq
/SnJTbXNFdO4d7ru1VgeqhdbCaK2X5ms+VvkrtxAZV3VU83rTtrPz/FcyuP4I7HH
eAfNeH/Rp/y0zrXCLvP0fYxkrqcILaidBdhIC75Gc8bXwye6BS9KvysDww/iEUOw
ziJN63xvAkZZuPbYMaHdr43YuupQgLo6TZufM5+KA3o8CaQgfmICB64IiVsk7cCl
ja3TDtWl2hTpODqfU8tYC21e0LzXpE1Rq75xBrPN0/zfMkeB2CS5U1t3zovQd+qw
+R5/4JWbylojjyUrLz+MXk99oITzrXkEj2pVEnNfvlFsOou0yPNOykYZowKBfe11
KTjHl0gcF1yg5XLF/M1pwqwAmdM7/yrCmxcbSvTrZz+W7vN7vTmDPPV5clwed9Yv
MoWvHlYU1Ny1mLynF+dGtwjjLjFLm/JfLsO4UTMGCRCzkfrxdbSHOFpCGcxMX5GZ
IWs0KM0As/qLIuomG+qQMpBjQOF6fnWpwj09mJPkU5aL4p2Jbqr6/kcAPIR3bug+
NqIRAVp63gZui2Esz3DGqW83ZqYHmykzsyeeJQbxZniopxagRcANG34nVzx7Ouli
g4LV6OLW6R46UoLRwXHpR/HJ1UVhU/i+q+YtiluPjILtf6uIvRIBDr/FB2ACTXwA
Udh9UXVe5slNoeuuZVGtxy1Xe3sHg8YXx/8evkYDLj28blvY/hSVhkhuoQZOFVj4
2OKHWijXMLW3+5iiI2LGgahFFKOPDHm0GgWTnJLl0p7xJ73/RTXA/Ko2oLzaaqCJ
3nV4F5E3ji4+Ge7NtSoT0P/dsLzueZLUcAJvYyrNe/4A8JtOCl7L1QCi4ZK3eGwQ
RblIc6s4o7oft5ro77RdbV0QHfBX5b732oBCPE607DPERQsSRulBE0fb01V5GI8V
/hYi/0Oynb8zAEGXySG4Wl1QlHJFQs7DTb/ggulWgYK6Qws35TWe8rSjFO/V1q3p
Ufc602NXWtVY8w4ap/yUcECNaQTO87NIWu0JxuCe8Afv6Y3eipIRSUo1JEEFiSHl
DfPa23hw1rS8M4C6QLNWVCoGrNLRVPjBElxWvVLlnJ02E5ZtyOkAoNv3AiVn5kc3
CkcdoBcALBPzw3oyGxGRzkdtfAGA77hp21g3DIfE/m8eTL/a7xcxitHDOza6qe1H
Lsqs+d4CYJx2y7EVXCMSBZxs/P5Hs1LwX6jdmhHUKmi9KGONbIKleLgujs7zfydH
d2JdAzZEAnP8smKi2WXjsfN7XGMR1JkU9rxXFevfGjNfGES4qw/cS4IkR8S9OsV9
+GoIMM0gvtHHcfTfqkWhP5vje48rkQG79RSOL+bWJRprgRNX3o2Ng7+Jf3oRGVTp
6Xmvn/UuOe4F5yAstWBY/FTsSQSR7Akzg4ajvAidV3jE4jwunne2oy5eV4kTI7q+
qMTl3424+NSRymVRhg77IBa3E2GpNoTsRwkpbEwxcrYucPAGACKGjyPvtWkzmA9b
lEesQyLFIPCrJqSW9KikS998T3+NT5H/4Aieal88z9nWcPqTaGgKxpSxy4AH9j6W
6KLc+BiA+7tiAXMcwYtlXRhxk6UAUoMw++OEkpohbvEn2GgxE0ZjNcIDSgqZ9X5E
uKOvnkiBX0RGsqflhxr3NUyyrVF0TsstpKOpkxDVgjb1FdJezcF40wEt+i7ryOq2
E1w1sXs62lJFd+jjtkr53QK+bJUZL9TcUZEy0G4ViG0Nr26EWD6dDpQbS6r1vDfY
SaE186JtjzEREUtfuMuubm7Hi21kWmQrFvg+Adj/56/Hc/Meajv0lQh8KpZ4hKWv
kc95gIKgMF1NiqNBCS6WsgSG41Hmo3+FJR77aymKCNkhVg3t0UTLOqAHYYLxoLJh
QyUwFPMiMm6PNHRASl1tdXS2HLn4jefx4Bjwf05wvxsifA3l9fbsq43YRuT6mgGC
mv0R806c8mIsEpHCG5qeHGGFjkrGQIA2OYQgQlhJRpbHR8zx+I63ilcm2RKDPUWs
OvIs5XHScw4CWulN+GkqX103WmhaerO36Q+M9UKj9aDj7A3KDLh42dioywc53n5g
ARfa9TX25PEDjDN0lVcy0YO23RKfqzj5rbWXYyy3GdEjSKNGqY6TxmsAgvIaG7uJ
cE8Ol9FxyviP3JKdFz/t/eAQkVkDKdLebfgFuZu3uT4pLYMTiW3pl6AUSdEpw6sE
l4cwFIAa94azQHdiro48JM3/6AezGuxzfQ1bBvTTHZ/Iga4zMZ+PjWwEMGBymvJp
RJvsKPvm22N6x6C0uIMX+QbcQ8a3ayJ0zWepehLRqsMM02H6/Koykni/qVTvRa8v
cHP2jaaJTQMRewVTZ6GGKqNURYBtbCK8JYpZZ7/TuK+26FRs/WdH2ovKJ1Iypq8m
DbwtKI7mNVai1V4CJ06wIL8Z9soJVhTpGedfS3Ia4OalPaGES1Uv9NNUjRHmijc2
M53L8zg0cPeMOAj3i9ArxXfcxl5UBODeLfft8XylOk4P10YyxyT6JLRej1/Jq/CI
EpqlNvOUe5dVdVL554DTkktiId7oUIBY+0XHoBTLK4TOwyMBEsYenxWjo/v41pAO
n0p0anfh1S5OUcHyzvDLAZ+ZIhpiLUlyFTcRBmX4Yp8eXefUoyhGtqTljsFk9lTj
D82Fy0oT+ePS4x7586RQbsI6fzuPVQdB3Hg2483RRM+FcaMSjkHSwmhJefF+UeF/
6dEWZYMpHuq6M/17ko5pKMuQAlCWaQAWlW0tw2/UtHjyOhA+3yghcYTMVLiOxzhB
sGrkUY8rRmu9WkrkRE1bdh7d0SxWg90H2iwA5Jg9BLdZKfabmFciBssebs24Z9VL
JV47pAbu8dR9kuHSh4dlunjFdoAb3MiB7lfWDSKnGkCcH292nPTWAqvlxX99yLX+
RTcDJ2gPImlSzVcJkrl3l7B9V6nQIUTGCi7gMBFB/aDyCZcyf9YHXmzfQB+EFsPp
LpvksCfH8TG2L9V8M1vpDQCr/OsZLyGat7URYPy24bzc/edEEIdhs352fZhFoEPC
zceJsmVquuXDL/HtYeUwlS991yRcoXQEtsXyyR3ybbhnFTFiTTLBX2Rds4tAB6g9
xKxQLRiFvNVa4oVtib2jgVN2ll3T6n09ScJ/IPBiDjjKb/2JnOxb6KBkyxEfUDTr
oeSJ1J7JpQnl5hGIei384Zq0NSC3PJQETiud5Wsri+jmwKNdNr2CWTOKbuMcpksw
VGubtEXa8bjh52lw10Kf0x/YtODhaTRjvevgBbixmt7/7yaAgY5ZVJQYBvJdtdsI
jk6IAnxCX4IZxeRQEQCB31BeGmsAAV+8Bk/xmkx6M4BBfKPX3NOcwglxKjdyi5lO
e2+rFYsBo6NOCtWV8yQGrpkzqzBfVcL240cGEMDB23iRyeBI22mr40FkpLYIzBpi
++bwv1+ZI4k6xcW/EZhE5fIkS5G7KmRU0NTlBnFcGJ+ssmmFAKtmQiLFzvKECS7y
/73SkDavXxxNNXdG+fKmRl9cmQfdnF/9HhDg/inq/GzMOUrutlFKQfXPznD/7b/8
68cNPwyPxelXuv18jkZmXH8m+PEgwGDsG/MPUg098dYmo0PPbH565Edr2GXzhnNj
H4f3P4RFE2pPY8beZffHmDtDkVoeaBO7WpABoMELM2rKDrTv0h0LznPlnvKmLK+n
VuISSGqQ+6R7YYpbsVxEhxjEmRSeetftBuRzMxlBpVsDPH0qpVz60Ryu0TISrCeq
BrilOEHH9KBXK8k6Csbj7tXlVfiA5BiSPpxvjXOyphxeg+g8o3ujYoArm/+e2XOH
ts3VB6L2p6K2le36shKTiO/a72Qik9NTNSjnnkTaNQ9qFfjBxXy6qnKQ8nd2J6kU
2HYyX8GyoCyJaismH8kN0B1f8R9D4rz0FtA04pLs8s6E3v0TKVTssPRTI5FiTYjE
zED33yJ3fh01kxRM03K2FBEHJFvitIrC4inJrtQ6P9tuLrEagtrkw1fSRRBci8tg
mvYbhK4GRHZq00MPCCoQkBna41qLc7FeMNnL00sOLV6LESbRC1ODZ8OSO+pujgQQ
X7JWCbJWLmDy7VzjLlzNSoN/eoICE3Rn0EUtyP6NtATf2aO6TfaeP3j11NF2c4Zv
jVgtWhF3sqjk2tnlz2UAl4dMfgHbh+rYhN6Q5TGMTT+ot/8KGgKuLg4jScHTVX+o
TOS14ziNLHdcAjD+sceeD6MRXffr5ykPsagCHzYbueWBSAIi2RnK0nw5HYQxOrFI
Y5bm2x9+EAZJRyl0yjvRUln1Ar3Je6P02+jh4jc7nu+ljOEq52EKTa8azxoAERXB
Tuj0qKeY8ptf5RWilm8rwWUpLH4LkNHcQJObXdxTifaESt5tfZaVoPQdHIBgoism
Jrg2ROxQrCv54Fe1qODfOyWSQAgo1DpVFPm8iwDGY50q32O7Qi0HOv56WAOJqXNM
73mLF3Z1kQ1zGcGxTOAB4JZNQHO9dxeXcxxFicwE+foGz1u/uvdOMf5jstLxAGxe
1gzEIr2uSOxWMGJrFVBH5OIBHDc7cn3ooHY3nLUSkqVmtNfRvHGldQ+xke3dC3gR
ODP+k16KOetU8C7NqwgqhsSj7Gh1WbQbz5gsq5rgY1VmmXgeFXpavcdenI4VRz/0
oFeIRm5Vgw2xq8fg8itv6pgwFVdni8d2Z+VWlvw0Q0SLUmAmXoYJHLQcuf+NnN/j
E5gG9XZo8mMPH9mWueQyzPS/GmCaYPNqjiYRLFQX9GNsmE7z/21ci8v++kfmLcNz
z/XSfhIld07L7X2O7RXaidHSV/dWFC0IQkhVKBluho5Yy/SPSkPy3G1AuOUY071I
6SaqccjvmUFRnUe3QrvdH1gclIfF9xx23VBLFj/DrDSuzVQYrb6c3sSWCCfN/Wnj
gljwQiS1F8Y4lfBnCMYVAEsa3f+1sWqX8SZX/in15HewcN/ngm0lUL8SjBCKRShg
eIZCE4k3yAkFE1FmGT09f+7fK86oUV3PcUk5jdvqW2ZJMkZKr7+6cuHzWnHCo2Mo
0BCeEVsmqdX6/zEo4RW4aBm4AxykFkIGXDeykk7koGiVydAA924c+Dyl0AksVSKY
Mfk4JRg2dgs6jRWBuYCY6XZ0QoFnUogTJ47LJSgY4aC0e6yypLU360JL4x6CARpF
HsApUdmOtdbAUWfdwpoKhQce7OmlqFSKnQD6FaXg06/WXmrZl4bEQLSXVNa4RtVf
fEQzLwM1tCUB0FOxE7ztevpMjpxoU1+eafbT5/L7A+D/+77ZU6a4r9BlPcZs/neY
SzrECVncvdJMrtcO+B6jnEITBDz9vbocCJP8VdETkRT/rX5m5giblJ5TFsUQ47nG
VLlhNAZSmqsIJMhVmJjCPZc7niH6fz4MvcPglRo8SMb0JAVJ1zj+m5jt+qq6EcCd
QqXXWftYPF7gkAN00mU5rbmdN2uYTL+3G/F/1sm5akNu4N82eM2r20ygSU1/4651
5kKB/ZuMRy+ufoC37GrqiEqVjcKJil6Vn5dMvQYzY9jBwRleJ6ySe6e4D8hM7tYv
U7i+UB4TROenqfZ4HNxneIQru0ZZI++Ut8yk4T/jbeLHagFRfF7yO/LN+OZV2JqM
Wvxk3rH+u8LFUKA77w3h3VgJZtQw2XyyAdpMj6UNcfJ8S5rld0YiuhDXgLmCkkdx
fGJOZySgQuRlADVivzVjC7Up9q6O3M00i0d6jqfVk9Pf89TCFQXxeet7jJ31u8gO
C3iYvqmVaZIkunZMRFnFt2icfkzBDkyVCBw587jvE8b+SGND6NFqXc6Hqv6pWw9J
8Z5U/1Vu7s/6reyQzUER2G0eiWpZtnaH3rkf1Hkx9Zfr6nZlCV30cgSuE63gOnJP
oxDLOwBPGTAQygXBeqmwDn3HJ181ZdPMfPinKfLcdDoD6NOJ2IjLhRMtWbLJ400T
31yDMGeKtGFTEWZTmQ92AlxknHUfWAhtgQNJBz2jI1FRCVqpThjrJ+Njyiplldnh
4XpuFvCIQHkT0i/71kfZDqrAjaBOnXjoeMzGs3TdNTCKSqnTSPwp0kaxelLSjo+v
TRaq2yIVptF7kQGXbx8C0vA4t7+OHdcEe501IJeF5Prikg864I3yGS9c58eGZcuw
MER5jlRYjvjbihX68IPMyNe7a8WdjwPO9AVt2JyN5Z8e+mYZOWoM2VrbI7OqWBY+
9CnbVp0+5/HgOCosFmx2tvuSfHR9VlfkFH0Cn6QmIJqdAtaZWWi8b1e2VdnFjQCA
GPsrFWwhMopdvPsd5g4Raw59ygj9RmFAi4oTNsx+TdO3YXdTtKrERePfoUA/1Www
qTX8ZMwqpntfi0etBXzTw/VUACaSJmuw4/7JofEypVY83b84UJzhnDgwYt0qZZVu
rrQ4Qw4ZdhnjC0gCSK8xyuSIht4F4Lwdnc8o0CzOngBnfxw0pSR/Zvz8LNEZfnAu
BLhxARfBijXz0a17NuRpxR6PLh0capkBc4O7NSYx7NcEl+r7AXBXOhpOoCmgHTnO
j3Tz24KT4ofzhKsTEGDN6f3FhczEJhfpIkPWdcngQoOY5vAJ70mH7zaueup0nToU
CIQWhtqNAP17gjPVcO/h1nVGNEL4UObycblFONQ3bKOwdkBA41Dw5ROMKBul+hkO
xeBeVeckJ6TxvWEVtU+8oOa95TJv0PlpFn1ddKFRoX8vgfGk6TjW/dNSFLg6lvx8
ip4IYZn6B20B/re1mA+cu2nszK08+h9WPwYgruSfHt09BLcfLqAzQOSI0G0Qj3wd
pTImdJEeniCerTZ7us89uuMz0zWJOqvDQoSlyeWtaPDzE3fhoKMGuVyXSb8kvENJ
AQoaDZcLW9OCDMxfGOW9Eu7+shvOXuhWN86ZJ3kwTbizgpxVhL5iDp9MRbBME21p
rDTXF+ojM+Qoed4AHmt4ZyBGU745/mQ7KmAgE6P59Tbbvqcr0B7Nks7l4G3/mHJc
sSGGCBd8Q1z9G57CmGvcBJ2jSSC+fnSTf4PQaK9lYLNt3yZ3NJTkjOgnlZGh3y5d
OdYEeA/Jgzfwg5FDhBlzXmhxl4DsKIl46AXelMaJnE8uzR4HRxJreVzbroJsyuia
b2BQCNTeILjhitqnJfvn75gQHNzRmGp9e9LDjYgy2vT+13PHdaVuV4f2g6FHbimH
s/9jH/vdt8/iqzB/l8Gwn0LZZZVg9pNZtiFCWQBFXY4JevK9aRu9mS0Smh1LRs9G
sGCs3wyb2Aa+Hfs+vNPquPwFYttPkul5NYHWeFhQTtWZ0EOfLme4rjFefE8mnvzj
lJKJ0UjPZ/2LenawTIDH4FuQPlhtU1Z2dxgppWq/2RupVH4i+g93+K9GXeyR0T3s
cd9XCoxaks8/hkZofwrWaKQLkn6HF9MoSK6XCgVn+HtFtwvOAe6xeTBzmrpusE4j
Mz9fSKEkxtjhU5YSUQJ8BvZZwtCsPtHzqMtgq+RRQkoK0ChAXukbhW/v+FoFIxmJ
0wKT1RIXWC8gaKDYSqToLfI5tZMfR4rBOLxFf0nUDwhqNC8CH3SF2llTjYBV4bJV
bWNZwcgAyrYGVPuKrJBUbh/Njadqifb0xc5V/tA0BIKrPbnO6vOVubTQX1lBFKN5
`protect end_protected
