module programcounter_assertions#(int N = 8)(
        input  logic        clk,
        input  logic        star,
        input  logic[N-1:0] addr,
        input  logic        JP,
        input  logic        JF,
        input  logic        Flag,
        output logic[N-1:0] PC
);

endmodule
