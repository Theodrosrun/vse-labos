`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Gl0GK/3DLDegCQbuenJIBeZHeYLOMmpZTG7fkDCjgN3md7APYB9hWkzhKUSSut1Y
k4+C3V9fPs6l4kBxGdxJbTJdlc6Z7nwHx8SOPEPoawOEKD7mpsgs/O/wsnjbGx4/
E5bFeXMCvqjj5fVfj4Vo6zGPCO3JCVQNOTyB1LQ5Qy9sY+tXMPs7eGOOjhyhdb7y
6TgB7iQ27qQEw1qNeeQt2QmNyaZKTkuc1PY4Jmng1vDIQRGdwW134yX0CKg3vSLd
iwVGjddY2PkXCdBtACW7ciehpNdeFbmRWPaXKQhplYMtDuA/9O6L1n16iEGLGZ+n
sk3VX0A81P8BAfbo5FQMaw==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5376 )
`protect data_block
UTQyfqGBmyxc32ZrcScnWsYoejWXlv3WKaIU5tDRUssbkMxHUhNKijCjM2l31qIN
yepPXQI7Hu05iRQor1ASNbJW2n/zb78Tc20B1GAPkokU6/5W7voagLyUmvzQw7YV
QBPS93ZUDlB5dMEyT4SpMbqTuN14xspNkLSvl/qKI9EP9cyyrA23K+0inXNYOrib
/Is26M7XOsGhQIhP+bPFX1vombvBdXQqtP/aJH73LCeLjpfBVe7Tyd1Vfj6BQfkQ
cjjg7s75L9iieS3pa0gC1sIArAOp2Nk5h8P+WnmZ7iP2AC5yJocE+/0MEAeIcuRZ
E3VfvuRozJuf8cXpaFIHuVqjUSJCysicnAuzroAYqMvkLjwsxQOcezb9IPDIYmGO
1GrJL/v8IrVi8LNWlQ+vLM4hszIwkAFC46ZFIgnB9Gc9dZbMKId+17FYN3csalRq
DrH7xhte3rS94yLT/RmlfuFf+zwQG1eyd1iMY4Sfhpbul4zIXoA2igHu1vS9oALF
cPzTnBAgHXbSIlSgGTrcOU6RQkqpbBTnHuzGj2cUCY9hMpS9DvGh3Ekvyd00jzKD
2NEt1kijQij29q17tSN2SIwSo2EqaZNZduK5Z9JuWPxA/ACCmYkal6OiLZDHW68N
gBa/V6a3gu+41mR3EY4C7i2XG4QTPI1pQ6eiLaBFZ97r8L/piwt2yh1lRCLZPr7x
nBMnQ6Dxm+1B8DB7NsRIELKfNmkI0TPFv0OMinDXN3c5L+lGB4CxXSZ8PRweabz8
FfIlZPdZgSs9YxMjUdmTAroRxoAEB+miXv5o4dFxYusoeep268fsSCoY5/iErJr7
YL+/baYkBu1RN/3MXFxcjMLipWvduhvuBXVKlwv8AYj2LeY82yYMix97Kr/WtsGh
kHYKlpBl18sx60LMt0kaqT9tXQhzFZxMrGM1Uqm6tEwEHIn7KmBausZj3lk43W6B
sMRwXi3gP2ptxCXgWOv/oKyqwP2qPamuUeaP9LwjBYF6wE08c5DWSfyKvTeoXF7e
kZAo/AzOa7gD6Zl1c0XjAHtfwab9AJ/x/Y2kZjl0InySnxxr6nBnxs/7eH7q14VW
Wu2PUU/thTVo6d02cWnv8Qr2ufMuFpgeHOosg/v0gJYLrAB99kTSwQ8vgm8MAlo5
yMsHK2blbpZkQGn9dVgFVI58020KNeJ+0MwGowqMjiti527gJtg/tmPKtjSRy7Sk
UeYtOK78X2xeIP15EwAT4251lqHlAHva13w8XCfeWLPMONdMwTuUEHkwuUB53sQq
HROFKaXPKWNKi0DedI24K7EXZULQZBMHh51w/dWt13VHIQAh8yKRDWmS1gTzULDs
I0fY3yntdiBBfOzqNe+WngCWXfMllPgZhm6nQ6ks6H29vXP1I0t2p0jBjYfons69
vVvVkH0zOP7r+I5KDwbGGdFwvLJM4qxkbgxUJXYEgxbYSt5vhuOCnI05jPyxUxu+
Dw650EcHrOrWEwzBNwJkHEryJbFKLTLXwTKcxd/4evBvFfYybQlPdQ+kfrLuuNsy
HaZJoHQrpxpVGak6PFcPQ9Huw9WAKdM8fXq1nngLsRIU39r903NMZAtAY3g7vNkZ
yJurGjrt1lQ3TsxsY8knAtGfqvlTRR7UDHV1g7TcHfOdQKdWyV1P6Rt7qhpC4O8G
tX3E9YL7REF0sx/wVeUG/ZRnWaZcgzrBs4mopY9dXG1bthb/Sd9M1NOno2PL682I
vLm1Q1RZHnYbEsIfyt/680yyA0T1w7WODbMPl+IktsD4OH3f88GnIPoOI5hp7sDv
RIwiFXGfwIqgzI/AqWsNUDCQK0numQE7t+terUrlvOL6gVsDhqStV9Zhtg5CoYYE
9yPSCCMz3AAMfuX6vdwXFONtfqJA43SKjA6W3TB3qE6tmaFIqkog7yXFQ4/3Enlb
T3He7ch8biMpx0jTM/moak7KdfzjRX70wncl9dVN/c8UEI3eebl26XjtIQxTHF21
ByXAl6Tg0CEfK50KVgp7Y1gdFGG2eRaiUdSNkoJ9fKLNLYkYhnzEy+nU2nObQNie
OLrEA2Kn6T22Y4q7dSRHhYdVIVbRr+2f8drYP9kIbdb43Bvy50sF1XcPuSM9ny/7
yzZKxOjaZvu2MIHY5dwf9u9uhCwo6PU31ZpnD2lLcfpZxXG4tcZ6i/4e9S53vHsa
J9pf3NE85XTX2sEQVRK5NDtCCd+48Vl3yUVItn/VGLzN0AxhLTLzU3j7sL5+R1WW
qTKpPckIsuInfP5P/mpy1XwNKEzVRKyEFnqORgw3s5zUw7VgoSh+xAw+wwFWDba0
+g33Cdm2nJQnME8jD/KJJhA4FvAec12+oVuk1ky25+/UQMyky4q7KZOoH+vtEQUn
YfPkOP7w04acPJxnmsMx64MUiqPB5kXIsBIJaf8bCN7O2cW+uotnsly+HfjxoCRK
+hY+eIXal4O6rS+ojCe/p++JegrVmv4TmzQyT8BGRE+IXtNYo+woooRsJVc21om+
dvwE6dDwD04rl47F0B1K7DUbTJyWpG6Uy1j0mcTraBQm8+rG7rDGDb/cCCWuV0PB
IjtHxR8JLRhrrtuKrMZjExwzSG04OojfdUKjphKDk1f+q6Wokqd6eANq1imIpad3
hh6/Le6dBUk9bzcESydtFHLijiAdTnBgWcWi5fg9t65XdNJ8DDMPKdmlY0k8bbWP
GYtCvjxcTM+C/NpDVuLqrDv1V7SRNdkTdEUb6EEOgtZgSHY45gGulG7h2Sr7LKdF
aT8rFX4zoHzGTLgFm6KyUrtx4ue+FVMkfcayJ2NCXVcE8lZxTBftzp35snI72i8Y
s99GfuNx8SgHFH7Q9AE37ymiS8S8oWMmCpmevsqPcn+JnN2Ve6CuT5KsvLJOkqIq
ecsZxE1gAzWJke0aDoFcj93smeOtCObjaPcCmLZUQpRfsHLCzJ9zdIDXpN5YE+Uj
RZmIqM4vQjeZOAOjy9+0kCW86t2K7SuPi2kqw+XdqOcvYo18In7AsOK1tYs/FayH
Xf2j/qSGqu7MkQZErNE9kidV3LmgFRLg463FQVyhUm74n8KvBu+zxAlkQp46HIL2
Xm3Tb2mM+aJjv6svn42mUshDcFyV3KFOZ3Z93jow1JAfywtiHUqhMFj3gV9j8dtg
EpNYW52wdMsAsdkpHpJaFgr5GhLGhxu+vxpI4OrYjT/tU6LfBAaHXMpj8N9fLdJR
sK0Y7L6HshvTlnEVaeKzHMK2w0BeMvrlVH2XghOhhst9nz2ExZSCUSvYn93Ovkww
UoErhG0ijgTtiM27dACAJqjULHvZm4OS+LmAvjirZ3hVZ4N486EM560KO1+KEWEQ
6NUjHBEYghqrWkIbemQVQOtgrYfLTVHH+H/UuwIRJdrffcXs6Dxc2ijxGrFS0pug
G7YtF7nJvNdUS8OplK00g9hsbS+6/kZph8nDVhoPqMAvu1HeLmmIJanCUuP5uRcy
TAX5bJLe6D1yHKrDRvPCTtxaYUFfV9a95AqN97GV+8ySKi6HDk0+r0iCyJ432dQ8
AdGuN+rqFEyTNLhtPyFXFll08ESjhkYgJevnK7k70hSH1BkzxXX9t792clcy0lLC
Z2aR1CcXmq6yHX+nPUh53Ldie4IXqKF3B/IkHasSc0xrbnNz2cVHKeMKIWOkNN6Z
p+W/53+/4DXBu+IpFABHaQsyb1xWym7uG+KdASOpE0cQqMGcW6Y9XfJnZzkuYrV+
BaWmdBY8Hcydv/C8Mzx369UAgFyLdUw/0106HRDd82Ef2D0cvp6WnbYHd+cV3yGk
GBU35BjOPNuOrcBkjnCZIfeZgVupE9ou6GMWggs0q/l6AKyY/OdFPtYiW1WEeYSR
2pSNf9zfQVEF35/ybiSOH4ggRuYRplXQF7mqvUvILOe9OsMXWhrzV3x6H3tQhIiU
jN70mEPtnxzKkmqJgIZTCHh2u5arb9WQBaGa0NaTX8V07s23YPQp80SdzprpRDUA
dWBB2SKAiC5A9IXxVOWJkFsi2XTwkSu3Q9Iq7XLvg0kA5ryxRAfILzClBv8qeFVh
m3PaYwwIJ+LOHivgZ3Ub75QyEpVZocy1CvHTVBVRHEZIs8fDJwVfF22yFDg9rAlU
FQ15loxsiYDILS+nMMI5dB8gDRPVQb5t6Ol8cCcy25Yhf4kPwxi1GFce9lXDdbvQ
7d3HsFXtBfSTBI0oQFPxGMKNv2xN3TYnbRuq0cTSdQvXIETtxov9qqzK3fbpNjN9
JlcX7d5q8RiBmy5WO5syYWGiq/m7l0TGysmUWSE+yGLtNLO/rB8i7JrkvdtNAnHy
6K7ZvupE6/BNQryum9B+0f2B9A0VSE2IEILxWCaM+b2aIhEf1uYeMxcHG0At6Gqo
cVells0ZnLG4ZOoVn9GlBCEj6QNhrVL9tJsvXyyu8Pe3oTmsSfbnCMCc3O4RQFva
c9sr0RO89QvT+w/NKnTJlrExvB6A9ItrNDJMgagn/wvvREKKOJHyUb5JQTz1t9V0
OR9kHepnqwDup7WgbSXexsha/fLleZN01wqeaGv5OJwgl/IC0ADevKJ8NH79v5Lh
EOfZMtOeSGxpEXnM0+ebXwu77wAO9SCT7ILzutuOunpEEezZ15DsuQd/qbl30sfl
yXhv1R/f6fB8auO8IyojkTVE1m4OKzbb8nkqEMcoMQKrQLAsfVifK99S0rOQ2tgq
RnZmZatNyjac2iwm9Qv5p0+u5FbiERPY+t6iG6VN4O4uGNU6N4jfe7rEXlMmBm0z
6OhxxS5D9z92vDXiGqYPIB/gm8wW1bFzdTiXxoiQvvfX3Y0d9Te83WLulfukmpmC
yFsdERsyarrv8NM/Ui/+jR5pvBbfG+irvDu5heGa43j3oQ3lP3/xK78+wqhMRyGL
ZqX1EPXuIn2LbWIfyVp8GUJO2Xm4LbCUIc65p5dyc2Ka0hDcPhTKeD181h40yajU
xGFVA+7fjNI2WhJciKfMFmVFywKUxxHDDarjh1nkxtOBZkEtZxPDZAkyZ/2DIDDQ
W0cT6EbtYyNiraY6B8OjRwLXEsIXczgKBjQD5quFzoVqOf0YUKvXsb1vTHRmTvz2
T/pZ+OdGAjhn4vSy5RESHJSdJHK7e2N7ndE09Zs26GT2m05kS52071LdvbsfCuua
phICrYKxJ8WE6rMRW1tstEKkZclPIJ4l/UCC1r14WOLijoZCmc3oUcIBP7bi0Hfq
GDm3/9J4v0lrHIvF2buNGxLvxrskLncrJZq+ZxVOx4sfaM+i4A/FYhpaqT6PH7Ww
rrfdMUAkLssniKXvw6/X43qOHCQJV4R1O+g6bmoTVkkqQLLu45Qu/CYCIcq4qHjI
elMM9KbWWyn2RCNxiZ153QeMJxviTN6h75C0mqVpu6Jub8/KPp3lQ6Qb8SKxohv4
kS0Te3GZuEEXnQE3dWSpndCsYtSg5bnlSwTTJVLxFE/kHvYAH9jsZ9P/iqiPw6JA
kirBYRinIp1XvKLF7cx+Q/PLtwa+f/UADApwMWW91X2JUyZaIR8UYOjy1Va7pC+/
Qfhz8hfpPGjG2tws0iZsekVG8MiYObfwTHvw814vDYADQlk1fJrU9dI7w12qDVp7
tmEcOmzdkLyrG/2Lp68eziYvQ4RBhRd2D9vgsqsGxnk6UVV20roiK/T59OINVh+c
0l9NrYjmdJMZ4/nJn8aSjksp0mdGCw8yN6a5D/1QUXPFLjOXvRcwi0SnGYOEEean
JxelYIW3yHlv8jistVPIBey3+Gcwssf2CX/Te1fEShs1tDyzgu4wBLuUECjSmwz+
zftAD1du7EaNg0aUyJtqpV4quAZIvlzAOSdilXS94DVcM2gyx5svJHBazJ3dJFUf
Hg9pfQ9g9Rh7BjS0r0GRQ1LzFra9Buf1uZRgORxTU2t9iskoBB3p3Tt7PSsI+Z6e
rBi9t4ubPCuV49n2ZzgdsIfu9YWnvR06oD7HWgy2G/4VhoWkHhgWufDuOy1N2QCr
RXKw3bcb3fbfs9LJKu3VV8o3X77vEz5pVx4OIkU2jmoIpDjTqtCgbt6ShDaxm1QJ
+yPllywLpXX7ct5fIzQol7cip2NT+H2GTZGqdkfQnKzMVSEyl3BU6x2p3DpMhynD
G0fYaiYT/TK13wWtVXIDiy1iuGzzZOJTAshtnD9W5kRG33gP8/sidFlv0sbOhqbE
ZaW2H159D5rWMfw4S88o5cE6A4I/Ef6ASok1r2AR3sOSClybK0RF5tMNeQWAwLiS
8sTjb6wae9jy9ZHv3xhbx+YpmdBJgnUs/x5ewg46Bbdq9IDgFJkS4sRgJkxG1hwt
s9ab6HoNmv21oGC0Z6HyKA8ruB3JrdfhS9qbNo+9uPvIokZv/qbzpce8hW8N28pv
KN6E44BLJ31Yy2cJ1quGSdLk/PRZ1BAb8ETLqM4Iv8syGJTVkT9kOaXq8Miy7zjT
xeYiLF1WLEbhzG10+ho1AJ8Iqyg4qYdlhyUWa1ZIMM3Gb8hnCMRfXrVC8T0ydWyv
wgL9CgcBfJBuPTwxBPZjqan8HWx4B5ox0crutIi8IeKFe/LdtWnno2lr7yXdvbxK
7u/nQqGmO+V899nwidkK2OdPS4krUTew2pey3AQjbSzyNv5LjbirdMMY0O33kOI3
v2xGKc6uxJnaRLIB+yuIRtRz9+zKLLh3EUz1VTRcFF1Mvptju9NxV+A8EB5N/YD5
ZtrzBe3G27r8Yz+C8zTXwWj9xHnChCGTxzyJZ10xsFVbq/ud38oJk/znpDH0KPNM
NJzJIO5Vj6HBr2GUK3v5A7CEtsUDk0RnvMqwoCCvR/9ob/JwiK/4eW/Rd6//1IZT
q17uhDxsRH4MDf0mpcYK7RS0w5WojXToYd+AjUP58pYLaaOAfSPyM+QvZS3CFHa6
sOrdswhtGJzf0Ek7L92k75RRsFIN19gW2AHHdO/sOG0LHfPJCLQeDmQSxinhML3h
7ji6eNHppsmPLJbTkD77iwgxeI0RjbM3dQSDB7ltK+9SOyo96M8JLjeIzt4DKXn4
njU+wi82KqAGlmMUzEAgiDEvf5A/BEd11yL/OvXDdchY3NarVkeKB20RWeN58aRh
SHtsikCOrOCsSJ5uuxQ60JrXkXfLs20ANJdD43dbKD5faGMI9q1LJmQwZxnRRjwT
vb38ZANDjTfVt3BGiYqRI6nLq5F7PyGlaBh2w0MbnK0ZGHxvyQoa1Oa17NtQKcyP
`protect end_protected
