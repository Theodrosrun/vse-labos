`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a4vAy0laBNnkfv45t8AQf73F+/ZtdvCtOqQ/MHo/VnWkPjStIqXQo7Ez0kG9xZrR
3oy067ljpt4c0YI2ECo27zh55G44Fv4lf0Mqn4QO89+3r8OUfdzfMceJVXDS0klo
ikwSGn+onNffPmGgoVVH+g8jE5Savh1CFAUrZIDbRS/5dNazNHPgPnMDfKLFvgx6
zaNGlEtEnJxWSetkAGtoZ/MYxWxrl1Qg0mLiVgwYQ8/kbHDvOXIF3OiiDIMHUla/
HLrnEihMi63/VGiK47svgGYGC4S2JcT74BYA1PAfvG5EbG6GcdaSpDRUqJEamwrx
3Wd8umN+UtELaWuFHm4Tyg==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10544 )
`protect data_block
2L6noR4TxxYzpwywnU79eCehyx9hb9IRDQOrl+7AVwfXCw0eq7KdKiwN3JtSzfcK
8TkeF0inoWAUMwnvrc2bRlCkna+7Brugp8cEQcYg3Dr6xn0qoGaQkVxKMHEyl9Jn
f7cx+kKk3P0BbYo2mqQGawKdCdtxlcVBMyrUFsMDnGnONGllq0wvKpx5o7LVQo1I
b40KHydntjzfmMBjt5VWGiK43TQRKYnov08j8bwl29IygusC6kNKsagwWZ448m35
ITbGzCYEDMFG4pJwXsp1/aF3HRbzFs5ak2Wf3HzCLAug8XmoNRS/6DX9YBkMn2ov
DdJrsHSmhm3SGEwI382mQvcujA+9a0RhHXU6d9L/QybqQOjFA3wKfPj9xM89wndk
jT6w3NZLPBesIDrHA8BNvW3bt1W8yUlmqU+47gYWQUkQK82wCyTXhz3HHRA6X4kr
zZ3yZTjyeQnbs3AMSdLdOZVj1xwuyvccn3lrcwQivax48L33toMLpvUdEbo+YwLi
p+LB62X2JgMsda4jyBViIDPYRWxLmCjf3HlcPu8YLqxiEtNUZtSBlu9JjUtLxynJ
U4O6E6EIq8WXqGshu5FcsWaUFntLJs4rSVWvhF5PfmPQpxwjhjAqubMMJ6OnOVtq
ipdJojkXBqjcRoM5pqThGBzsuJYKwn4V/IDcRpKqjx1tiqdwaQh22gadFY3NH/OK
XYTbOp8fGCiJsrPf1g+vYkmzS5dgaqx5vTBowTRZIMGAssi5a4mS/AabSc10k7ae
qbtGWu+Yj6rOJN20NP7n3iMd9o8UKXPb54iMZ4wqby/89YV+snyMl7g4eDt60rpM
0gV995MctmXDO/SihFVkeAiQenfn5tAnl0i2FK2W8mPFv1+c2uSNg/rRHKQPlXFr
TWXBV5euyWlpFTKAgaKTsaBml46UULzuf0bHllryLcvFlHqQbolHmQM7H5XL3bco
BJPlvBX81WbPZX+FZ7xXFbtRs/UYbV1gOkkyRMTVS3QQ0XR6GXLChPWfiEp77hX1
8PPgu7lvFdwoh8ZQQW9L9tdVbwc9BnfbEC3f5IOi/70vmHJ+1HjseuMzzb5QVFGq
m4HgYKNd85ADoIvgP2w/nSDuX0P9Z6pqS6QPwGtNwJofoyNpYt/zQBbj24TGadke
iEbwnp0xWDfWSH2OOdt4pG5XMXoT/MaGL3pvO8sP6XxtOI0B53YtjE4xQtoYvlz8
m9XsyiQCPvp7J3u89x2kWiQEP+HF4Z9yT1uXPkbcTXYQ8Q3YEYuhrYiwUzoleXUw
99h0N3HctNr4BIarxletuFkZolUG2TTAvPSi5KZdK4RAfu7maiJH7beNlA7hYJUJ
lshylzPIpN4kF4tlKRix4W2kwuQ+QqMZ3BlbH51CcZ+a52rWJ/NUm12Giki5xdhr
xGFVK06KrqBB3f6aON1XU3fyNHAEg7HAXkkWQlUQ2wWx4d2D0ycd5jOOc0Fiw3Jr
xzuhuAyUUox43cWeiHLese+QkBP6ZnK+pc0+VMj5nhNvu2g8Dg4vpAhdNt0M94JE
sD4EtR9GjJNx3WFOltwWTdXV2czg0eyUMUVrjA7VvET4eGhGWx7UPQsEUBfZEHxY
eh77kP4WbY7veD3bH5PCfrA1ipqUlgXxymPJwkm+GnSp1AHPFxTuApkDwySaBygD
up4+O3hSdQM7wMo/1Oh1ySE5utm+LkhrzeK9KsTlO1JR18z+MD5snITovbb4dlBO
JAU4dS1W6xF+E/KoBFJNmqaQ5sEoH2wMzaZ6K5MZhGih4F52eVfylEoQBjSrcv22
fxK6jhCr4YT/Bg7JV9bOAZpdPl4Gw+no7qKoIdJgDzKtEnMZy1h3ecAgGaGUJX4F
/vlBStMIhj+IE60C9+MLpvOVqdEMXbGVCK76K0dNCVfvjs1PnBqO8gHUOqh5fLUb
OMmYrntCMRl00dJoJNrXjhDmN63XbWGX/LVW/Aa/kaHdy9Butkx7ssqVdu1AVUYL
K6NflZQ50wx/TLq083AfsdEGhxdgXH5UvJO4palHV2zBFXzKBaRziOY1J/9VKN/X
AS89utbUElkIU8VYcoHMq5/zCGRWmYGjfYhNexT3alfldE8rpYWpKvhQeFciDpdl
qjOi8jPWCYZkJk3lvAiOh2/LGzdq8jxeQQ+HdJ7T4j+J3aaBkHqyifEtKg++SMJ8
x8zKtgRkQOEC6qRev2MMBX0ASKF0JlPzcfRbPUl4Y7/tqhSyu1FI4ep0R6GyP5cC
PHnCma5A3U6t+RsZxWklMwxKi6tVAk5So5Xyd25JbfAIe8vOBHc70/ukWvbDaJXo
QnHrtFAeOkOmT+fiLDK5dCybe9BDr9sYjHXGtoqEutq0tn8/xCzKXEWF89eXHchg
rw2EFI1iFbUtWb+u7TbFJ+RNeK+gqKF6JLXD17B/ncRwj386p133XPF5DDBCISpd
WHV+6wNeMQgPJYElAzy2As3zSumZk8BHmNoX7HXslmfhrMwlsM6iRWCBqo2x1rx7
h4/wv72Eb5WJl2lblfRd1ikz+sKaYD5cVvbs0d2au0I16yP8BqNsAGMe4uo70fjC
Nenm5jAE8A35Mpt4xgi4n44EEzV6cswh8s+KnS/fkICIJrPg9hAE9Xe3JRc0is5q
nLCZDutsEveV9Bx9M/RZtg+26ToZorEOMSDHac5MnEaCIOmoc4xQyv0WymOaPmph
3TGw1P39CTJtJIb36T3hD3xSupW6VMne4qRPSg2lzf7vbXrOU7/+zAix6xnB/sKD
04v8SH6H0h3p5HRjRGopxleRTDwOU4GW29tBUYHqVQxF7wljAPxPh+hPIrUPuhmi
5DpxgMPH38sFsbGX52fZe2EKfphdFdZdjKGIkq1yCqiXWfnmdISYc1UbQa+8ARgd
ltR4GMlGm+3a2veN3tTF/HHPLR7KnPRXfd4vYr8FN8X8R/KjAQf+Tj8kqcWJ2OKa
YFTzYN3xttgjt5FSAX/lE+5b/cyjjb4eqKB66B3LRwvuFcpiXLOY2JFYzMXlgOHa
W8oQhomqVOx074Ns+AtKpizSLWHDg5RfFa4Ce+K5DJimtGqFEFYxBSp7WxMWd1gG
iuTte6Oe8XQ0RHECk+rvMFq75Nok27oesIx5hcFPAKB/Geaoqka5HW6V8HjQHjPu
v7paIFhsDfk864zFCBKrZpeZp+xGwFXwxtdOoX/kUeBKO2CaSMy54Z1oWPOrT6Ok
lzqHHVMxylBffPtPbBLO9HW+0zV1r5Mj5JuMChZkPsvoAWgCgrX5caNosuyZ+IR9
EFk2ZxAViGGo14zgCgTj1/0CIrNhZWl99pUdtg4wh9OQeCXfJHvnmkSijnWogtvR
48Bi1sK3kyErsavwwjzD08y8H/o9aPvADWZtxtSsJwmyDlUMTcioamNu7VKPRdKQ
8J0gstuSlP7CImfx8eyMD0kf9BL42Mw/vXGXttstxlwB9aPM3/54AThUQ/vZ5GAC
Z0cEDdQtMKeOkcka5gCk8m6SFfuBFuWqQItjvy4ySppnQCYGP1q33mpFBCdi18Kc
Hjluo3VtNq8sIvYYHu6REJITjtTDI+mB1Klw2NEORuD6Tr/iwxKIWCUli8qhTqD2
CcFIfXu5yTK4mJczKHYZaYj3zXo96jRZR9M1d2YR6TllDWP1JkvfOrgM3PgEshEf
J0kgor2/bLhLCJCusO/iDN/Swg/A/5SkriGtVvaVAoKNU1/R2LAekqlEDf24vc2S
yu4htXoacmBXuJv+zsp5i4x+VLb6+d5uu1BwWVSbilXL06BLq9mdoNAjBYirnzXt
UpXlMUUVx7xnAypU+KaUrfvRXNPdfKFQ5aTk6mqu0aJ05tvN+cIvxOmlQmeiE3IG
gHpRWCcYFSC4vj44xMDIlKGrOIGN6BikxmehoBwVAHoCy2B+XpRmM30gMD2U8NVX
mi20hRq/V8YJF51z8c963LRBkWrhx/rnt4wh7XeNXJNmaD+uIEWBUMCEo8Knv+rQ
zxXLfBdBz2U69ieWorNarRM2z0s6LAgG4ogZBmRTQ43t6TLm1FawYEnE6H5Sdzvu
9nmwmub6BKZ0bGhXv35GHtKFGrJ4NylREYovXc4AFTLiUZi72Sh+0FnhpT9vLpNl
8bNJEeHVGTbF3E45l+KoXIUA0OLFvgb5EReUUunIqfauStivWFXq2j7aelcjUDa5
U+/4NVs/eARJXa98JJFGh8rO5EUBIvBGIUmJ7rZOoUMVCSMyX0Wr1JxrZbEKSLY9
o02cZZjjUVM7eD9G18ghM/TZMsBQ1OqQZyTEaloWp2OlS/vRbbL8ajRO4hVOjlzr
mOOTzJmy4G5sPEOnvK+f4OK6dEizKSkvIL1Ficju939Fc7O2sFxBSr/uv4sc1DWi
rMZHCpKrREqCMEmdqJQFVlxqeNgiF2AFGYX7EhFHe+XNBcsz6FM/YInVLzwYbzSj
6KjL2G+ON5RwL7lfoVmkP2iWT8rEHnmK+r0t2i2PeqRZ3oAJtzpcA2FnlKwPrLRh
jFmC6TsuIlsQ3LHblCPy2CCRmEf5fIuauCBG9eD0YSQmM1OwVweq/VwTEgAf52aq
te1AxUblU659Q4cRdcxzTeLmse/rtK33MKWEkVMAWRF/mEgM/KoWcY7rwHGL/ecx
dBG2+lldO62pNMaRIQdfPTamGcQqYhUkDv5llun/RlKcuk28EoAUMFfg0fpp1LtP
RIXGTL6II5WQ/vnxeu8s+Aqon2ZxbAaag19uNu7hHly8TBKsDEIvZDd9zqkWOfF/
gVzhmrD8uzZ4eirUplW/Pp+1oEm3q2FEAhlatSZ/U9Ql7VK5w/XAHc4GkLnBnAKJ
1wxgpyUQmevH1isZDORZ/dD8KPugfFwpT0cXntUXgur/OpW82vhBptscCitsOBxo
97HLz7qFkbM25WJhwdby8LtM3wTDWNGxtQO3BKPmum0hYJxMTIEKJfF8bUqGKV0f
vuDBekeNzCimJnPeK94CVoHlDsQjVeb7jERl1guKb7cNxuDUdsJOauCkxaKfoROt
A8TB3WEqCA8Fgm3jRRuYGRTGo6u604bAwY6JnhWSjpRVEb/kLzApMxw9nI6Uy5SS
usl6PjwdcejaML6/nNNHy9LSblFZly7bHTV3qnaBaQfAGhiVoIlX+hfsbhGnlSzC
IZ43XOplgAAk9dHTlJ92+R43KGGbHyb5Nyyz2wiFZDUN0T5P0ByZD8kL7bvk7h5k
4b7avtJjJUPF/TmjvxIIqS7I3bTsGmdVMIP3cuaAyKhZTBXkkPdGtHVDsWBM1oGP
J+GYdathLepRNFJ/1I9oF7QxGGFM0EeG2u/ZLwsw9E2K4wo58onWBlv6hg/EYTs+
Ymqj1gP5gekEx3VXwtovW7702tqNy6dayrWxvCeYz+zV/RhYPeTPF3XsyQ7FNKWy
S+xQyKNRGeAg5Zua43jVa5IHqVuVPT0tdcpVlkdiPsZ6WcSXHU+NA9bCzR+9xbp3
UTe/L5YWHK7cYCFc7/dwHuDdwev15/Zg8+3zGr+F95Q2EyJmKJiqPmRA+CCHm0Mt
bG8wIvjXQaS+T8ztoNrraHyljd2OlwNoNpsHpmjTgIAcO7AJjtR90xCo3n4J7f4J
c9XB6DF2cKQ+CQ+F2FaI8NuIImsM3FUVqm7IJBonyrXcrHeKcwbKolrVgB2vXdL1
IXLyiuucoBwjCzjE2F6ZVnNs5/fIAqfWOPhIMnpfl1s9BPEYz2burS2cR0qghrV5
2vSgv90sHu8ZGovcxUGqfM+SQduiKIjRS6sg7SyCF74d45+donk/1pdpwT5Zhzv4
Wm3VZmJK2i9FCS6Cmy5+gdt95rmCz4MdVjmm3fHOK9W2777dSPljvLE4BxKMKmJ4
HNsEJtcMbUe0R/Sdp9hzXCj2p8YUfvURzdTlX+fBqFf3efhGv7oCDEJWBlmknVwn
vVrRx0t2kvczKQbcjWx0Jb/bx0u5ZkYeewA5PHXDCiu6OkQJNM7bjoKmHCDTw9/v
BHeCfcc6A4R6kNqVETHkD6WYW8V6BSnyRf0rNnJizqmBmbhiTC+SQsFdD2CuBAue
mIcRrkL3v9dMTPtlc8y98T98Dc9CfPsEk0QazZTdklpA9PD+k2GJPRkTxks95Zi4
Fn+DFx/B6Rca67jZz8+Qc24Nnft4glvtNfR8frCxMgFjcLF2cYAIruL8ivHPdvp0
aZwvHHOPdsM9iQIQsbJeNAQ7LL5XgYI6sfLHb99ZJzhI74g5EspASW8LKzpxVHCf
RVK2EpRgTQBeBiZcibqIySG3i16Qdtz3tXLfvB69t6sTpHCwtGE69OQlodYsntEz
cw+6blvoxEk93cYWBYhR8zsYP1Lwxbye+LZ6FG80DUBsngBXiBeqm/hbAAA2sueH
leFozB8vCp08WcSnuqA6g8GHGrQHqVdoiFeidu4KwpKr8uZWjISx046PaCaO6QON
Twc+ZFA36toRRNQY4u5hooN8Lq+VMuizacJEoGLPvFO2PRDwdFHsEy77lXBYG8Ac
qclkNuUmBpeTpl8soTbJcbXK/+Au7OO5CsrnsrJsGNNCpiUzth5CI82gxMwCgpm/
drng4ruwO1LkyJ1IyX9ia6XoL7sa3oo0Y5Zs7vneVu1U8kYgyzjSGzjREwiKw8tv
VpAdxALmRR9keWvB9E5p8HL8Xv3ZuHASLy231hxjoilATHQ6EeCTUU2uFGyDeqYZ
2JzAUBw3zrx3ol+CIII8ozX5FNnqNagWgK4r3ayg4VAIcqE2donC+1Ja1zwkPTOS
04X7CLhSmYvfFViJwJmBnizG+MesKpqckaMGfU5muqEDRD9wkZPt9HQt/gHZHHhG
QUUumel6vmWguLxYMfRAHbhNY0+kbmvTCjStQf7qVU7xhaWVs+q6hPnZIcxAlVJo
Dtm5gUePDaGekg3G9+aKHhFxsWyiWt9JVIJs7uGaj7XQLnCDiyAL54Ftg8oTFcqT
bkftXq6ueEvjm+CtVePaWH4hAFTwOu+Koy6UVmWcg1GpA3z2ltOdxLjxMUrwAc49
91xzkNuB2teJuxATKTdSZnU7VI4O/r/6HRxdaZ5xiLxiPA/ye90DPjCZw4RFU7hN
HQFNJ5YOs6t/+bt0y+yHsGWiVEQYSoFZW1xLVHk3hld8Hh/1lip3VC5ww+Y4q4tX
mmfUEBAbJKPmXZtImhB9liXQVjIIF4MVRS4eUbCTfqpCDawVy1fUxCNlvSfm9fnn
RrpVCDeVA1YpgQ3M2Wef+8NRw7W4XmmiHRrn5icsszkYstyW2S0tYlM6J7AU0Vh3
9ADeZ6G0/7ovDxHrFVu+GfiMW54hjWPmSmMYEY/yoXXMXl3DgBn9zkgYSqrNn3gI
ajLmrxF7r1QpucnO0UP/CraEF8GL/kNIy6Xox3DtfJn8CRB8w0OdErcc+8EeXmgk
FYKCBNRqPdjLLCFw+vR1PZrJ5uIb4ZWdhnEckvlnlmAN979sVUEU0ACQ1PTdKN6e
h5723ahsSXk1Lx9XTG/j8h+SymYhYaEmPm1bZLK26ElXl986t5PJgULbmiasRpe0
OJH47YfTYRuGPWEWlrbNNVG+wTXxScICObKJOMWaPnUkdQ/UdohHvc9ki54Q81P0
rDcJm6DCdNK4WYqp6f6tENPsV6/+p1fQX1qm/6WC8xNI7e4ibTdlJzpp4UA1gBk9
Wbrgp7V+XGzBzWyK0VQZr2hA41NE/1EhupPcnuIssddTfhAfPi0vD6vqXKQLHYz7
G7bBgpAVRy3mQT7WzfzKkV47T4C7pkygtB43CgSsvNDoJfoDLMDyJnrGroNOdy+w
trgDjzEwnzpdxJGYjcAcbQNQWUis4ZPnF/9vSlCWXLbxcpoyHex8hQWKPgDF9oys
6sIPT9rwhGmqdqggyUT1SLBIFWd1SGjg4DfE8WcguA4yjkYd2UJs3K2MJyJ93THl
jDwQxhaFMo1c5wGZbDEZWywVE4L9tM3ch+oh6FNwpL3VdysHcP9YyuBaybW5EiOP
SuY8viR13R/JeNaKTceLd8z6l4LCDhpzgGotJeiCjJNEcteeGNLEWAy519itWj3N
/w4PRv9BCtVxxmVwAiJmliB+5pv5uyXXTFIxvEhE5dpvPRI/raT6M93Vf4GRNGxm
Z4Ub7I8AcvxG2lBbaQjpB1PYxgGqvAhnQHqkiN4mue3DZ3HbXd/PcigYtok3fC3x
WlNzraBMeeb9UxTclxWZxt8WwQv5uZHIXxPE4Yu8gRWIX5GXC2kNdfdvg6l/CD6W
mAZY1aHe/qhkPh8UvNrmWS6nkIeiW21pbQwFNkoKj4gnj7r8dP4L+4yc6PwLPbJc
lFqWCeTZmYrCwiCSEUYinHHcqeM1kCh693a046esNtrPe87j6OAZYMAtM6rh9Y1V
3YilnZzafsCk8juZBlfGS95WI48W0ORVGAkg3rQFxz9H7NHO/0/KADSK8qI6x19s
aMYmX6SH/NkknqKUPAPPQiFMogAatOLYZXAsah/xOlp/u8F+qAps40uE3CrHgVCU
RpuaNjfPKZKC0vb3ozQznYPOpaOWtq9TH/N+ytmW8IVk+Ap6nWa0j+QG33yEItHA
xyn9w0pwkqvoRgVWk3y+yxqnqnJdaGy3fhGwYRbq3135coxHATUgghshO5i65225
6CJDT4TTALgi/lb0QBPCxFDq2JT/P6XavpMGYzei24XJm7dRmvMmmtX6crzUbAgc
b4J2T3oQRBeRDiibh4yB1INzg/3iSTyyog0tMR3skI6i9t/r4hxthhipLTnnVtVZ
SDL7UJ3L0+1DtHUMAs0cf11SjZQ/hiGpItaPpLZEwtePNuRhZ7W2B6g+XzRkZE8z
cO2dxFr+YXRBMMTx41L3ttO4/ED7X+WWVpn2Q+oQb++n3nBgf38YXXoipTgaMueT
heOyYDq+xOjshRDiYv2C3ffhRAkGSbfWN5i/eDGXWaXLSUowLaq+Z2YCbXrtA/C3
FCtE9kNz1Hb6L3iCOsVDHX1LQ/vJP1dA3rIs2terE6CDOfaiaPMAopEkR/VDHwiz
g/w996NTnWdhV1U8Y76DddXT1VJc9+5lqVAwmBkRAhp8V6shsg9xoeHBHkVsDyS6
FDopu+Srk+qSruZCrPp4UI/j38G2Zd4wxA4nEMesc4MhuoXHplD1uT9ITIPOzQFo
Kxo5QpD4mXsfTZR7w44N0l9UouFu0g1m0QkfCTD5ju1qPrUaJk+sLzzAwVHnhZam
2HG4Derz9RSMaM3hS95kT3S8tHcnaxCWDFlfLw+XrjamqY6skCMFcMMGs0zc7i+H
bRv43ucJHTQ64wUJQcmhmDKii6vEf7sFVHILRkCrmG01ge1I0HPyUYukkjz8dx4T
8hCnvegOc2KcD6yTdUnQhd9cHqQTymvCVHLqJ5ir7/Z3SukywzLWoqKfUBHlAkUF
Hdlg0oSWCJvV2pmjKp9jsu177Vcqq/fCMClIoDd/BAM9gs4LpL+lC6HtwANDxq9j
SthPLgQ//eUSdiY4duDLuFkpnHFLLexCLwPiHdKXjb/WHPe+O1PSo6CIHJOxS9CV
dC739nkW+pyRSEbmBJWDfvK8nc+TIuOqMbJNzgY9iGE3LVssBT8yhacw6vcNwE+J
A0WVN8pqhqOEC1GnWtwo4/2/YyX/mYLDP9KffuirrUloohSCK+bl5hkDaDS7x8u/
OwY3tvR+UHNoOlSpqnqZiIzZp8/o8cjiFfC3gx0X+DuTSDx4+Gd13PGJjHmPUfEM
LPIBswFoNHZApcQh9p5ttKRI0nHJWE+xvbmzWPcbK7uzQ744Sy+D4OoPGuP7iHGw
ZcgGXsSK86gc79OUw2LQjDMSyBbNUZCBQ42cOvBxU+z8xvWLinbpH3LKfOQ3rgKs
8FY4xzcdBMYquAjJG+rYyehpI8FAIgD7o8s4lE1NqQcGOVlhvFyAlDVwchqTeQ+4
WrB3NHTFMyS810sF0lsH8qSOdMTIVa+VNn8aLGYCuTXUpgVh3dK/4YeJUpq69rdA
QBVjFvfUysJ5D3KCPpDMr75ctVvmRoXLyAvyLbncm7RrMG81LBUiEOyQFXLfqXK1
405y95WShS5Q6FdrV4skF7f1RLcvPrGZUek6DcUseCjUJY0GaEzVnyjKcFnEMA4V
Nxpv0qu+5pEDoY3cMF9k4Gdm9AIJN58a28bdM+7ZKWUyeP/XWfc6uO+jEzTBamrI
q0KoKpCPD0Pn4XSP5rz7AiJWnwGpaqWMfC1CBf823bQcaU+TTJ78VG9pFrY2LUZi
VMO4SQJHBtUqn33BYKJKKeZKiqYUPzvYslxXswB8j79zYIsxbvQ6nu9ELEJzHty/
a59m1Vygn2yrczI9eOi2ARTV91NzL5PlCsDUG59RIVIyAzDDDL00iBRqO0bOsgHL
RaIzqBKHvN9ce0Tbd294rE6e4//kE1wsx5kq7JBdeHanSGKLpESfAGhf8aAfhT7t
KL3YKQrEHOyU+3uU0fr5fF9RhdXwgkk2WR1x3HpdWh4PGa/2jovYntawTShx+pDT
/U0lQXDsF31j8KFc75Uyo04/6w6no3mQhfaP4iZRdAEabHRQhDl+3MU7y+pg0uo/
0K1xhAydwCVp/o+JI11eUZ/bKtacue7l6R2lKrv7v3OdaOZ21xFbXAswGXQjJ1FC
z8JoIO9dvOn6GwxFTz5k3J4KppbnbKDs0BZ6fcg+ez27XV0o05lqaVEZFBg66wO9
Vomg6UtNgysUam2gZpL2oFOZrMtu/WQt1cofKzP/COoTJzDzEz94bUJwNyg0DSHH
CvmxgDTvw/DHEZXSp+BZvICyp4AdR/xZlOdFBR+BaFKB+/D2+DMh7cFK+pPYRuOr
ZYgvvOTcNUVDmtMO5RRYmYxag/+Tv9V8JNJxLmYUBH9AfvDdWwuXOvi5aaJyKpSl
S+KcHAd0oeEWXHmcCA3HpDi3HGA0vkr+vzlHES94t/3AXbGaO32WM2dRuc4lUguS
HIaRyGa7lPxB2O8g91Z4dJRpN65tG9DWCUXJ8m0PRj1A/pQcM5E0oXqBhx7cO1cH
ZlHt2GX4IQknOhRkV1g1EOwcWzDtanDLRgjJt84MGhP5NBRgjhll5NxUIVW5A6Yx
cPYkqHUk09rRiqLnSOsg+Fmfn4jkopGSy+r4LsOo5dLJqc3Drrf/DizVN2QpnKqJ
E8723K1TxJGw1eNWQbk3O8NaQESj+sd+gOoFutvVmbeXuwzFQBfBaKPcO2kgB90x
FTPmxfjCWuRpVbB/w2lzp4M9muQeBo3HOcO4Krzfx4IxS9vABDf5VqN9DO4vwn8y
s1/nOo6r+OlubFOAl1In+SmAsSjgHj9p9OykwWg/yHuDh/m05sqGGciSSRBxBYHh
lIlapE5xrbZV2W7bzy3O2VlRCohN6NCPGjcYWutd9PZWSEykHNTz9Ty0oA65ObUy
MZeIoalTFySxsmrrsjsuRlL8fHjPJ0XriqsC+Z16lHkgenABgRONM+8SuQnSILuP
5ErBa2gEzTwtDln/eIlYFAGgSiTvcHhkkpdLTbRUKfjfdV+N9BqDuPxK3dS8DDg+
qPgxtpw6yC+D38a8MH8Y+DEp1wRbLKXo62qiPl31dRxyJbsmrzpOYyRfG6aV9dbs
/UYROgo8EMIzFUpsBwNjVDKWr/3oL83ZGKNlNVLsVdu+jU2SR0On8oA69Hj8KTur
MzL0O6/5Ap3fJAed+vjzVwygx5yhN6u9FKbRhQk8pXFNij8xus2o5EgpHh4TzSOi
+I/QcdxJsyty3s3vCiKKFqNNZB5qcxP46Men4sxmmDL0wRda+8kt/UWOzKYFl88s
z5MhHG1I3ZCTO7B5xmUMkqu+3u+jHB9HRWV0BvKHPYwto3KMkCIZw7PN0CrZ1V+5
zaWgD08GVGooD+1ky2QMo5VN04bi855MmW+rn6/+x6ooXBJKzJLx5tPyjLBiLxtO
RG0SGhmcPuduqSvEhcRe7m/tm9o0iujcJKLQrklZ+hndq8vC8yC+LyzKLKYs6zSg
rLhOFsCX+Fxfdg1djKrDzsWfrL5+Y87kGPNJf2cv7enTzCKXPr31Rot0bzUPBm1d
GJhmhpzihSVv027ysTYpDRyWdLeb384S3hv9TV+/x70VKgQw0nQ4yFIIO53TnmGk
q5Ts2IcZvJJj3xZJVIbXIxEQETvmLBEEnwN33JKRecaYOdv7t/UbzOj3subOqY57
1Z/IAPVsyYtJy71YtSZVakD5HPcXH3KO9XIVw20x3HHqtvG2KgEt80OXSvBOCmM6
WPRx4FaaLyxSkjE7qlA8vTYbA36lvlt5rFdEl6vgF0dqeRYh2znxCZ/SXlIz69Jj
Hpj+Gy29mjK7lVR4f8DSyoVLnC86cDRm8zEjcuS8xjtqMD3QPa5EqfXKKW/AAwGt
U1N15IjNIY95RHmYybXVm6fLWkSY+jbwWE5nMIymRgkI4GT/YwjAQgYFSJc7ZDO+
TCnm/Ni7vfaYKiJFoRblrohuOgaGbD7WyL2Xjq8TLB1R1NXZwQoIr337MGT587i4
QRNG5GJ6OLcFXtSC/VPUeG7+9y1KLwp+kFNTjTJAw+07R55xNNwSDVd1Lobrg7A6
7+VshM5aT2VpWGyl4zcuOs8KijJU7CJ7WxUQ9Jb7Wif9w9LcfNZAylGmEFFCF3Ze
7n7bsEeOptgv4TCKRh7V/Lkqx/lw9v/wXQDaHLPVzy4H96GBY9Dd4r5XYZLyC9T3
48V5KkcUHn/8PF+kWQ4DSDDLcoEW7I/RJGHpA2LPwUA3vmbzeABhCqAM9ccPq8fu
quUWdJxGOXmsWkJ22FtgItvBzv71sEFU9/PnZJoFssLWWpcKW3uTxj623do8SKqn
h4RlIyG9Bc4Dx9V2TPthxU4/3tK3bptbF+kEs3O6AoOkV7PdWywXFggg6BU9VLA4
48urJVFRja1H+HG6zHnGIXYdNo6bkFosa5kk4xBomAlDGtvalOrcSKGnWe3e9gYq
l1fONDxDaHe9ZCVcGQ5Xn7jlqaG67a7Fym8XPfzEwOk1MO2OeNr/44Ii0dPaO+9o
qxb4heKXjyDKwm3pKsFzO1NUi6qvyXxAq/dQz8wKw6xvp8A+a9TenjoASwEScRQp
7CaMUUQmCfm5NWTxW+bvid+CwCbHgmlWsoF2PrIUTC8+TLooBBnnq5XUeYrjiMs3
/Uk40VCoK9J0uXbjsCBPLcscEJR59c+DE3McSqnT/Ar0RjfPgZp9/7BFRdmZAbnA
Ysqqg2pOlLrvbpQj9SixV/oDhEc3NINdxgVGgiTPeYvHJTlQ3m6uXgkzc1X2EPmI
nyBa6WIrcs0GNS8Bh7yaWkDLDIVxh+JZhEVYuoWQm0hnFFI/SxHqggqOElBPrk8o
u2aZTvwAv02OJq5TWcett5gEg3sH7fBcAgOFWg1KCKyDFW6TVbEyv5nSjdTG50WK
XOxIgxBa6fQ9qZAKMWgWUZRVGc3HrF76anYJeFvUZI9k9ObzG8sNVniv11ZS2AwT
B2Z5VE/sCJYyZI7GFVr0UIesuHXkoSsfIxRGAjmTBGmtrd0pGETFZ73HSMRCVp/N
1Xz475WzFvRqt4WTPNEnP9hvIno6diR/1ZB7ecunSPdfdl26v0AiKfdei1EbrlhV
MEpM7w/DJ1J9cBSIIaThnQN2w90zomx+9gqnMkEIPNF+J8NXbqbLe3fmkjzDoltJ
CB7Dosp69OZgSGv7c7ir9thDun33uqesUal1/3t5q2AA9XqgBiQZ6aUApSIq6mV+
HLehH+AjP2yI/FI3WD15EpNOQC/DTdw1UOB+eNhGPnI0Z2EO5syVXSdUeWYwtPl4
XwX+LeHMv1evsRqXsKqHIV8gCBs7M9oqVJt3htCA3C2LHp9JIte7h/w4XHbHFMIY
nUW1JjyVbMH3YB1A2LwZU01WBR4pmjTMqv+kGzsBC0hrXxGAczz5kmpiNE6MaqCu
mK+F0ZCGg1RwvA0lan8sRNbpNuI8/IKdHAg4K6Fzj2X3BjMcgyOwziQ3TgF5+YcD
lZg0p+kiAzkgNQwEKGZxfpsI6YF312WQCpSEBB3peF+GHRRcgEW8bi4qbZgP32KY
fdQc5QpFkkywrhuZoXH3uZ8kXwx1zT0Bc0G/s5UHhDK5IXGkc3/YrDZ6UvJwJ5NX
hOf3BNlFHODvTPw/Ke6XjIVb9Yq3ZyHREJu0jVjDWNQ=
`protect end_protected
