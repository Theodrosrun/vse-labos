`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ADETXHTQ+KII49ZnXDA5AV6DqGXNGD8BYcCweY0KDy43ONgMZeIuf7C+PaiFNSNx
c/8R4rHTeKCdbXbdZXOvU9p0BPClhrmpLrGJehGBkUs8BK6GB9wGEUAtvPtoutkY
qBiZi7siudGbjVOil07XixVjiTVioTX8k1sOYBwNFw4K13GL+sy3QY/Vr6iCb63u
6u5W0AIP6Z+FMXJytbUSGCQ4ZVUsm6nTcK3XXTmeViDoVZR6Os3EoVj4VTw47uK1
IwIUfSWlWqq5cue5jt81ov3A+xxi3hTpHLCp/pCvRVkUvyuIx61CUo7ZExj9ybGW
kpuZbnnsxzhtW6bedApM1Q==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 19136 )
`protect data_block
HZb3V+zhNxb26+W7QCo1miAgqA8+zvAkbZFrzyq5TZP/ootJ7UVwnmlT8k5y6PHo
MLEcskHJhbkVkr3OyV0Bx8N599IMLmmDGFcQJ34K7AQQbsFbYIegb6SJwzv46bHQ
Jb71WeCwaAN0dPMTgby8d2ZNEmacSH4aWvKkJYGYR1LDH8Jm69A67sUbbOWUyd/8
LBrYHEmO/6VNyA9xZlOMiD8VUf1FfR/2fTk2GhC6RxY27qMCCY0NP62VjlSFXRYM
i7E0LV88gkzj5Fmtkx0jT90SdYkzKl19vmNVCkZ1NneDJS7j/vyJec46q7kZ02o0
9jhR8Gg7IkFuM/63SktjtJ+pV1ir6ioz5tBFtXEsZ8uIfqn2b9Dlyqg7MdzxdQGH
krULZxrJ6Z7FU+5SnC8LtnlRYZbD9OZrm8UWSEZeO344UTHoWTeM26Z2ZyCN+CiO
T4ijxzJr3OdQNk3AQg8wM4C9mxwacGXTu79AXe0sbiH/bZJTnF1v5fp4D5ATFxlA
UnJWy8iPuPRrwuyWn86/5MXYJpc5tgBaZvpOUS+5/H5W/Ilibg/pKyfvkgawLOMH
0P341r4v7N5agbRooj8Dx3VlxE9PkeMidubIzg69iYW5bXqN1FiHQ4TCeSltPc/P
fMdjOJbXjQkHaWXBHDW1fs0YT74uaU+kuTSqP1uaDW+yHLOZBXjziVgjYCtCHHB6
4GayG6m7O/ZhgtJfUjMIdLGGVrHcbrsGn0cD0Ch6z0a88PNEjVXTGYg4JR2NzWLd
Yc09c8GIw0hXneaSoydBqzeJ8WBxm4TGy7Ro92G/JmT6cKjPPkecfGCCRYaM+s/s
VBRxOvARDDJxWwKZXne7MwrrHcyUU2m5Ta7AA+UethWGHMIxnfrO/yICRjkFckfw
pRo3DvMdVAYHUlfG0a7Qgta1OqsYSeb3fBkU+aKm3Vcl28N2Y+TP3a9S9PeVcPTl
RPSZS3GwFwMNN67cw+peITDn6JqXjZ9bmvmmFKWvMkoAsqs1OBy93dyPaC13EfV3
tR7yRebulgcdE322qlqwUlySrcJvTLrf8aAgq7tK4+6ueSTjcF39RN01FZK4BRp7
FVyZ/L1OyLrUXD0JgSI0bhwfwoIzh4Km/KVXR9vL589Pbu8Ow2+ozMiSyqKTBcOD
56r/wPMGonBfmgXEecwFCRKgzIPVgzrOkTwc5qpJcLn/gI0m/UVhJYQJZBxrgS+/
Hb3jo1ACbCygFKlhakHmwiwRIOQ3kJPkKgJI0GX+bG/QtFt/0l6XUnlC+tJ+mCiO
VQNFJaYm6Qufe0efCuFBjD6Ew3QNkqhnPAjNfEiSPCDwKyvu91WflRaX1hgryR8o
wKeGnotZeEgvQXlbZIR07gRXhUJ+B8Ne9V4l2VkXbwHGIl0PzjSABy/cHjUHmR67
MxLRTByamSWlJ81+5uBSEveRwHpgFC1tymb3UX8A3q38AXEojFwdP+4O0SIeo2/W
CVmwWUpNYMEx5ts3GALsyWxIn8ofJvsncB/tgqfXg+5A3Iw1jVko1z1B3Y5EEV7I
dVS9/MDwHKNbq/lMFN6Jjaseoxhb1yIOA6TS05PBgUW+3xdnXbuy6g7KdRnAQYTW
Gy+nCDu0hr0siyXiliK+EjG5rtShpeSx0E9fUcED68zICapwvB4wP+VXefUcs0p6
NBUwK10tr9DQlFn610m4kqSviJdd8f8aR7DA81ldlW+zC6UdlhG/60hU8PQtA8AN
6mVpBjkHmHea0XuUSGCYRrTZVIDJMAfSWhMTmAqF3eLO6bK3vRDZEaolvm2VXLVP
EkHPe3pv0+1TJU6ZH/Dbe0sxvuJXJEFCKMqZ89zKMbfSu26EPmwpuEqLMBIBfKDe
b9JG/jcd3KE4TEQNvJenSt+ajDhbkuV6IYaXodn5/NnLIuHa+1joHwB0EpuZyxde
4poembLAE2HgZqKwI+RalqOVY3GP4I7ACgRJdYLB22hjV8FPIxrYrk0wtHRfwKsL
1s4lm8wCdB/DqCmiSo9Ed44rfn/wCxWiYC0QYuMyMqafGLs4Q38ktvSQIgdmpaqb
T1j/OfEAp42nyb0+17qxQPWw8Gsoj51zB2sxZ6iqqDwtSpIjOF5d+7AEuNte9xDs
wM5nIR5rsW/JZxJr6MunSQLKnveuTUSgE7qpzRKJpJJGdqozIaiBzjT48NDx3P+h
SNoxcPNOnUsxmkTMeGZqFTg6xF5BPdIdQnKfuJh0PRbmOKRrr+idjfURUcpoP7Sd
h+9vV3hu8gVHxhaaLJetjN3dcLnMvnIHJlBzbhqWttaDrvqCm9uwHUbEqDckAprM
USbBsGQif5cS3+9uJj7i8IEUyQiEcK4y8lE5CijegvW+ewIV68+uzE117s3Aw5+x
yXR2zlJUHnulXt8drLgTwdwyR3/GPG572iTSNoB0e7gAQqf/Us+CLv4mVcD9XH0A
+B9fvQ3r9tDRO/+uaqLQDY0mxC2IPAmz7Bgb9x+/ynbHC/gVumzqd72aV/ssynya
KtQaLCh2tt/V5pemr+uB0k986g/h6eHREA6NbugdqoRw8fJM4rZEAhyvmYyZ0lsC
sexRmyw+Zz/CyAE8/Z2A/O89EJc9cm8e1MUODzD/LxjE1KqJk+saU3vNW4N4H8UO
mAm0xQVpzgE4I3+k8UuP38OodE+0PEhdGD66ejL8tfEt990H6Wvpn9ZZW4UirZUs
0oa90gxOkoE+IeWdPbbJ8/MnxdsNc40Q6ikEQbXs20G3lMGqaGDLkW/3pk8TOhkk
XDEL1A0tfCccOGSrv901CYSU6ePutIav7rtu9va2iKd9z98K/xEkA+bGFhyDQfDq
+ecYL3Gmn+9P3W/n30oBk1zuDhdVKB20izNx8ub4ff10wrMLAFU3W4WMfvYE0pVO
taqoa1V0h3AC7QU9WMiltEdpJq2hY7yqBM0YY64H7UlBLgcPz4R54Ap1eEtkf6N/
FhyEP6nOwOPzINxTfAP4PHczmfYInvo5z2DzwPP28Szklg86Z1y2M07eosUS9nFT
DJWQ6Vd/PFq7SIWHi+CGXkdIPRMFiBhS5NZMhE09Ruq1Mlmqm5NTa5ocu5vEuENl
tI0HfGILw5iqJDWcr3wbBnCZUdzbZCtKBJvvhc1/aEjx9IOQtOhDdUvfsFYRvGbq
5X0G/VdGHHIeqgKhSlLm+qB8FXgTjqpx24MUoKQuruyhoGPPVO7Kvt56O4dwGPIx
KTrdq3DY5kS1Wv8OdWcfHSVvJz5xWIme2Qu8giak3NqkMvjS3U7kHldVhJPi97yA
6dJFxpHpnPUmfNo7pnIe0CkwnVnwuk1CX5Ms/opgzHJC5yNZ2CQ1f/7sbCgGfKpk
MWna1sVVmn5U66fHuDOPHsLSK530FrDecw3apdRdItAQw4Z0f/nSP1VkA6dgFEka
AskqjxtX+z6ylSFawO43lDd4sEnDLj/GgzLJisujwRAszBYdl0p0Tkr7WobfB+RC
ryEee361bPYygtR8i3Ucckkx3FDibAaWhQOH/tLOyGoM4kdeizdbiKPYRsAAdn6g
La0MiWuEODMRTTgxauOWOLDQAnuc2kNgpDEft6wZTAO3/Q2bVf9BjUG8/VZz4cEj
kGfgLcH+lmU1VMTeJYuVWQ23+zPzBoFqzk1hiteK6rDlew+bqjcuwPNLw5tE2MLD
R0TmQ1ct8QuhurFtIx3eRj07wqBLcLcJPyymd3rPxiUYvdtzx8EmnHXRY9wZf5jW
8fg06DdKXD4uQX0HcDCb9UwbNOFdMHnmNea/GHspf8m6kfG1jR8quOyUdQBJIjyS
rwys8TQNP/opbmSr0sNyv2rHL6T9GffGtV7m5IaGp3O7GyySGL52nVMTjQEUzUyf
jZqHuD3Mv6RcWJkjbj0m8WXBNnfgJOKxYebwMqdAJKvFL/y/bbR1ZrVa69pHWFNo
k5fp1iq9elba67BQcz69PxKoSaz3o22jVDzOy7m4IM3N358pChcbOoWc/z/O1wF8
wNMwuJefdOXBXsQTave9sQIp3VfpPvArrBhVrYli62d/ja3PiyX2sokloYlffM/q
rZvUBg9fBP/E8L0Q01/1qnHEQ+Vbiqq8zkvKP3haS3ViZorGmjZN4l6OAtpJKLPT
LEEyJBKwpJHC/X8oQ2o5RxkfJMIVeuXJrpdrRxiBsUyS59E6Ovryuiah3MDTo+4X
LMXyD4utHS8rVkbUA31kVZVAIE1CBZbHaHR5b7VZbcJgsZVKAB2zzoLRKQG0UcIG
OBAIDpyrc3kqoRNR1sBqPSvGd862T/gGRyCP81sVBD3pDMF/WboLL2bHcs+0Y0kB
PZNhZEt1xlnkxpU4RfP3yfFyQ0hUoKVVfj807rKKnJuTCJqk3OWqwsgeuGvR+rYf
FoLoxSLunXaKgFgZHK7dWRULlowmzWGJWSatzCPV+IUR0L6ERp2Lvpuqr9bfgJOG
UcJ6p+Ar5vLh0q4KsgxrYsIiSaC1lj6QC8rukd+dTqFCcM41SW9JwVokcm3EnIer
tmBbB+TjSpyl/aiPExfV3V5zfHmKDhvWZ5KL9cNLObYxyszcbuFfMNQH82y7Q3k4
+YB7dZQI36SiL6+5EfKTwmHM6RNEey2ONgE/HqLLcheJoz7goTrj0uz+OmE/9uu7
t+BG17SxtM8oxVHDnsrOmYvrx5ABNVpzI0vocYThJwLP6nYpyqBh95+Jpj05WNP+
jFI3NXw/mjll+fGoOO8f9iXBgnSGhQZX1IRM2KgCA1Jo4/CDo5+4xFQAKAZChA8E
lJvtiJ/3tO7eCnzUZofpyjkvdePCmnKislTzVbnJBmWwmuy0fy+Gu0rb67YV+i41
MfkpplMq8Rgml5qUDI78MH9nUbNlpteH4+jwi0BRXLBLneYnZH6kKULyttGpHevN
EtODGYSkCcgUR4nPlhxCfOocVrXeCbN3y1UWNMwwYlj5RCP/GZdd/i8qLDjfvjCm
a6oGocsSyB1V9l+wuzVzSlCmQkctqZnryl1jrgFG/6uofsRaBU6EbiEYafjBCkwa
fGkN4GadcSB1CITJ92/mr/RXn4yQBjtETUIJRLbu0/16LlOhum+0dqAl0Y5eZovQ
gXwAhhysdUe3zH6JJ1uJxZcpIQ0WWC6Me4Fe4p3gK3MiYYnXbpRHDv9Soqtg/QyW
7BbfkjBWhNAMwkI96LCVS+ECBDxNfeWEEcYzctBO0bE+MEafOFsnkBSsN21gB//M
yZ/7jt41cYWtkR1TE6X4frgZrOe/M0y5w2yY1jkm2UP82v63+BRHblV92hySdy+h
XlLxe6xyZkcJZ+4x5bedMYXXbOx80t+Ewfbvn3t+8y6vSLRXR4E5fJk6vF2RaHBb
URXIZxnkHQhrR2qQSw5pn5i+9WepKblbnKK+L7e6FvuHh8Q8SvafCVYPCaQOgXfa
PpPu62+YnSHjrASY8ya+/UXOpG1SUk9bL3fAuxR7ws7eA0Zyc0m/a3I4Ch2Z2jqH
/O8C99GPyE/hVYfOhTApKltA9tNUsNK4OIf9vkq1QX8l20NoWYNJA5OrmXao+9cl
XC9W+GSbTAxvt8TSjpDXCbpq+TJCk6qVpSmS9UYFXF9iAqf2DOWtmvkJfx3g1C1Y
HGpNraPbZ8mgyQZ4V8vYQ3igIXuXk12tu7Uyfy7+C9Ir8eFluF3k8CRU7O4Jb+Qm
rPPzvHnYJplFhoGfBx5GGUe8cTmvKT/3Mboih8gtbb9sxjCvSl0wIZgu5jezBu34
fiIJoQjYVsH707XyKm4D22p5xI/wESXI47VhTqJ/pk2YR+0Ugm0REucT9Uw2f2ZY
L8Mc1KkyK2sPVDokKWfT0VYIqvHHvjJ13/n2QP+cmV0+vGPw0GXNdtroSQrHpdA1
akEoaVQusfw7oLD7iNjaS0ye5jJZgMUZuEadWUHXk+8XASyJlvC5OAoMJcs5/+eY
kiYVlJhe9OGCMFEcsq8Eor1+LRY8apNqIaj1E+eQZvN6xmDv0K+QVRAz1y5NHH1V
yKpUDy7w5PCuKxOe+vh+Vo4+yYk/w7RlfrhWoM0kj4n9SXnVnM4HY2cxsKVmr6Gu
9xUN9yhcBNDc3o6GvW9EBqSzupGgrVCrGToquiuzTQkAuucP4EgqInge/QXjYjjB
Pja/SAuHV/5vrJrnDawuQYf47kIr4pUBXF3Q87OO81hTlvZAiHn2pb0yfaPQErRf
bQ0E4APDIkklvHiwvTEofaMi4BeL7RGtWpGDbi5/RKpzpx3MajACodyxp7tz654x
cKFaqJ8neoKiK1o1Q8meC4+b7d9fGkubuXBfKcgJaFE/BGJKxZcvdysSQgzy7yjo
2ikatff5tVOHi21pPrbpn3TZocgFTSGCDgxT9bALXPDtgtE6Hr8wAT+LFfWxyFv7
g3Ypt38KedP/mtDJYHvxKVLFyRJMLhz2IoJz2zjIUOusqOHvlO5uEOnBkWXEhhbQ
NZ6TTs4wT0ISjnwj+EO3/o5wQhcDmrPGakV+6eeDOPfnn0LiMZMMiFfbEtACw5Yg
G44YcQmn41qk4CVVlttYKpcP0P11i/z+TKYxja8CJprZVhJnwBvr6sCyPBJWSbhq
0h/7sMvIu+jv0dzTCh3g9vy1AbczeFs99Bh7G0pcksee//xXr0zH2ackKicmpfn7
bgdlg24jCmuYv+r3p0LVTxVvZ69TIxR4l2JxNaRpcynnocNf5ym8jy5fpzc0/ITC
+VruRtOfX0lF5+Pfq7r7C5ivEyelBfCuYSGMVsYqRS4VagpCTyFo+A6xc16LDF1d
Jcr5BwPWniUgefGRYVuVJM2HpfJxlQB+O8it+g6PBYvUmnWAzXZ3zmplCkG711JL
SSIvYUT9LCo2Q3V5ow7fNe76ICtqQSTozOZtgQ8mD9s95luOcHvhatXwllpWm7cl
D7YV6Xrcq9pCHZ36RJ2WujJXY27NCUDWhsRmv0sgmCTnoCEo2EL+pOEvwNzUXNKP
J8SIfRy09TOyrtb2eKc5dwNAKILEN34tyWdVekA9vKhdvuY27l34qQBxMi5mcKaK
cNBv5KkeGrP01TmcOW7wLtPAMZ/PRuPLCrKbEkE4ZyCFFiCGDZhFzaY+pyvAwVTo
yFessLeWw+SyQ19o+kJBFTsdniESsFSFNrvzPVRyFREDBGwEICfuXukeOcNKrHyA
R/xmXgnibgi8EC2Ee8JHfvySrSSwgIdH7LPTl51y7HuI0KuvCirvfF5Ql9Zmmlae
DtkNK0vHKx4WQ9mD453/QRf5xndx053I82ZbdQOXKjda99HziATcgKLnanB4H/G3
eWZiUeZrc0itzEKSlxZks65sfsushEoRd/YrwvvgY97EuL0FVRZzU4hOUAfIYniG
4EtX80f1J09dfRZc4WjBd6CZBZHaBdGTDGnXJDmhganB/yDmYEFe+GOQgG3MNCHL
4teYIUo91+d+MCsIYUh8mklxFqtAES205y0Llk4Op6xj9FWtNCd+mr1Aysulchb0
UlPaA2qUPPJsz36QKAtjyHAO/rM+6iDbrWKhrTj5yj2tFRwVRQqpE8BT37ozYA0f
Nj9gafjwCFLu34ZKrFlaxRnXtjg7f+h/AhqL5tY2GqXxay13IRgOXof8C9TicM8S
iO+sY9bW12djJuN+CVMAKQvCpDibD6mE7/HKYqLWMZVwbWa8++QCitRsZFaO0ilr
LbcmOebefXvdqXILPLoC1e4n3xxPsW7sYGXklod/vR8Zh3SRRx4L3s8DbXC5LRfi
v9xBHRhx3AF9A1qKp3iNwv+AyHXvXNvVCn+ABu/h38fQGUMzqmz3K0BVui4DDuct
F2PVftB5g3AiWksJIEK5LDVPJsYeJsMU/K41WZwieU5POgdsS4xX7RKkRJRyRDxh
6hixggCXco0jdNDedxKmZnLYyfZIXGHfVTJNdQfd51kQIMevwiYGz/2xiaJbSjY2
Ux4LhIpQDaw/LSogqU3myfIA5EbUfBPXwJIeTc50psCAZtNQDJDGt2elK+TZu8KO
kUk+noLmCASHGTe8YlBBsqzGj9xqAcyw8IkUunsrJwGiIvhfGZ12icjS4MhpANGO
mrBKoeDtpBumzf3PjcZ5WAci7q1Eujq+GgHkbt9qPIpH2P2zMNWTu683myLr1YAi
TJ29ejg4R+4LU5R9zOxgOmZiVGSkx//Kyf3QkD4CMKkuf8RyC6a/9m8quxVLG8Ue
+3cNd8shAGGGRSh8iGmPH97kUNxWMbzm5wT+9JG+WDfFFdbNpR+ZhTLB2Ub2clZS
IQAzXSoh7vRGdEBRXNDbtbU8wmPQ8BHWGab8iuhTZ5fwlFye+AU0lbflSgxdGgPs
T/Pb+deXVjKMwwex5NERfD/zXuZ3qqHjq8x34POFvQZBN/7QCKWSGbGSatpeQHU5
psJ5OWquT6HnqBoBIsBvGeWHCqUMg8DTwtj4Iqg2G2JyzJq7T3+/5cAgwcH6TwSZ
0FiEDuSPJvCasQKibBrSBU+MM2UlCG12xVXXHp9p95M+soKxcMFCvtFJxKhiCTWh
goYykMln0q6kCvDGlyE+OxFtPAU7GwQCsEntaLY04IwGAc7KRGTJo9uHGZ2/iYIr
e7MYsDexiqRW8WmKfNTKsQhJoV+JOi5KIPmAR+rzkTzYyCGcm9FAaYzFGBdyGLYb
X1k+OtFHDw/fL0l352kY7J/nqmTych8yaKxYy62Klb7z8cHAzuP8tuTo4HgHEGla
L/z6WAodBH7fNxND5pIPglydLZLNd/90kybq3OSs7Y6eJIS8IquANioA0W0+TRzr
MPEb0CvUy2OKS1GZYm6igscBMYiWsPl4mYyQCE3wPU5b7xeVHojBGPlTYwB7abNa
sNL7f11LBWyV3n0biKNV/Lvoi5TH7jRfwsqGfd9rK0YslFzQgEBrW9u8iYMX25xP
BRA4UpEYSfvCNUf6ZvPXOpVNHlt06UMuqUxSlc7k8AegBlyzSoxGfH1KyIMMAcQR
LYWpWNafxooRxim77Xpmru0G8MAeKSPwJ4/GOIdCsof42ydOZ0B0rxjnYP3G0oOC
Z/5oiYYI0fbZE15021lD/FCIEDZQ7UrajWI+StMF9oVffLEZJHyaxrMfpH8vbHBo
pV1t8bgZhkBSQBIpZizD40n80E+GXeZOnkXrYtTJrpzYNGUgTswTFIGbQTMI4Gei
Jl4eVx/RGRAjzFbJR1uTaNVBt2T1Nw7WRgTdFrlN8K+88tTDmaAbmG2kFyNJWp/b
dOOYobdc/rrCyKjztP08rg9F4qTOK5Pv6rGHEJ4JvyPkny3ff0yVmA+fXIWbw9gB
t2FjvIBWh8IT6ZEa/uBYR7FI+mmgJag8Rae1UmpK8fdzvqBnG5qoV+PB82gYNf91
shQVuXKl+OjC7W3FLi+W7hMWvLHqUKGD5XYeg4N+Kvb3M6/fb3PyHJ+WWdNaAKUN
9xwgZb0UfcE3/KJN7u9xIFU6wZ6buRGtLcZYtOTVbLFRPvSMXSKyzozmCt+ToRIh
c4HVsBnLZ+BcAlQVfyiNBw0jeytVZvcHndDKKUMTlA63E3rEGxm1q0BBK3Gpu/V7
3zDviF22A/NyjGRdjlE024guy0btTydxF8Qs6WomI62oGC3/TUgpQbz8K+onOxsv
+mVCkf5iQKyAU1WK/wFNSzS1Ytucapuxi9x5HzlNOyTi6r65r9fx2SDL2eOn75ib
XKZNiKjoxQFBTfepdQnhOYHD3wz6oNOit+2xOkZpuj+oFUxKAI5WteiZzAHjMa/4
nA02s0a/QvdkDt0nUF6ItvzmDeX7ub0HSUnRY/q2X4BbmJMu5u11uygGAwHo2WZ4
g4K/2hR083ab0pncrEtdZijK4PSJe93zXQzvpwAuMPPLv7jowEwpCmCKikMhm9Jo
6TYYhN2ArwZxhrfVuFXXHYBxkF0QctkV7xNhdOn6Zh+j3of9tpW6IrdmbvAwk5Ls
OmfwxDNPwFwVKv1UYZDGjUXE3JjyvzL57HR2+hLleX6V2czEZTzm6fMbI6cjflY0
bHxGjWK9pRq/LT64aASjc85EgVm++3PNt0MLHZN1u3bKtSOVLckrLpiDF+8WKiRW
yPWSQ4fam1DS90ja64eb4rDqs4FSRdklr9WFqZkkbwYI5iwJarLZtEppDSNJMunY
Fr11ylqJoqH36TcDAXuELpC+aq0w2NIxLBVfJ++v/9u90MPQxwXPgOoY7pCpXAqW
phWdSdv5PoAg4QlytrMb5UBWZ3UnDXBDywfHdZ5QhR3XaV2waEopsVn8HV9x2Iwi
xvehLh+x4TT9Cd1VmWc6p8zt+Uwxx1xtnZ49elpgEQ6ULDwIMirQC8S3yZxsmCf7
VonlW8Lki1PSSJTZ4jyZPvf+9CbOTNVzoiGOU1nNaY6gOgCvRTqDfusU6VShFSoX
v1Q00FIc5s6w+cYlSuFgvmEvAzDr0rg+uOxez5hJrVtjGmzS478j/xRPhu9akvJT
Vv3qmaoOG2U1h9OHWInS7Jj0M9XP59/omlPrxn5XPM0ZziPOJfm4rSSOs+A+HP5E
W2XwRaHnxP0gqee2FfeXCGt8eUBPTfhgNS5I8FrVjJgmpq2MRbbV1SpKVifNMNCD
82RRzCVs0MutQl9wOZgYZG9D4FZ5n09OeJqRI9TnYcQhifm/O14T1ec4AQ8JvIQO
6uyAOdAm5IwLUqC/X8XHSDRZsurZLsewKzyCfIL+BU5lcLIOpAaM0tUJG+/z/fO4
BJNPqd+ChlyWQBIXfa/4DenoWddEsDtMJZgueHzAFmLizdVRs+5ad2DOFbKNeg+8
7g0hE9Y2a8aSNxGoYIr6TsMdWELKGQkE4fo4G03tZas6PDmtqFUhKGRXwJsxjbOU
1F0U3wb0CDTA4Li7AsqT91Smnzbm/4f+4ipJuP9ASc4ERYv7CANU7XewW1CdPPqQ
M59wf3MF7wYAwHn5kJGnHJTmUmVZxtVPM8veYnT0OAPGvWhBt3mCOfDlLhYOxcJ2
IJhTBWmJtNygTpGPY7zJGVYzcVqyIro8S2u85zVHndwJV86Z504tGaJ60D5g+SwE
Oh+vcKwRLZJkj5m1KaqvomQa3+p7Kt0Tqv9Igheb9kR+75jSTYreg3YPbr25Rj+D
SNSdhTmmXtjVwbeqBIp2wJIx0FrT0NSJMlBzAC3T/iBXpTrt7fgkDFoZjNF78a2S
x+1mCC2z1PvkjN9EvH3HreT1fe0JoPzyoUaXK9EiXmrePc8e9LLoLWoKAa+gBR20
bQAHHswA5DUDL4AdQnz872F39j3VeJqppORaUEiWTz4Q0US7UHuZ92zm0lfVUB1z
GqiEJpmWxZGeUsJAkzjgCt/3fohsSaPmYE/kp5plE+Xpz0mZTkKSzPeJguIoSqex
0ILEURBCaVHu4hh5U1jPJ7VkvAXiAEe4jPpgEGhZN5yI0XYACAPMrcYRZUreWc60
cA+6d9W1CdF/fFQJIMIWDK3C5lI4kmO0UTlZKoXYmicULlNLeLYMRzoqHRz6963S
JlcpsQysOnOGDnMADbQb5sv8hdLR7OGv8uHq5gSLqPwTIj6mZ5jHqf2d6vrvJlov
CEYa50Q/ZsNCMEVKCbqv26s4SECc78bw/gCtwRmiC5WX0ccgNFV3uCIAByoQnbol
GU2u/49WNDMKZjs0H8KMYXmJJ/4NTjgGg+5DW02hdMeQs8cStIxzOHRW2Q5Dozwl
7EbVyFEffndTpvh55C0UK4DLxE9k5+li6T0d+cohiCEW47+uq2nM5BRyZjvunyYf
c9iecM8oHc14VKzH9y8DWEXmqHEiWaAht2rAIPovZZ+kuX1bPdEoWCL1KdW4FoJ0
g++7uq8p0mSHekKXhVM8Q1vMBb2HgFfECvpe1nSM2KpttW2TOO7fXsPFKvZJCI6/
YjfcIH2b+tg5tBfF1hYqqgwDRZVDbtcnMC75INg4/83oKupXmBqJz6D5/Bg81ZXA
3nEn99aQe+6jhlwvwTiKTUnDDHpD5JfT8IJlMhWMp7VcPhUurg5U2PThK5XGk92J
VfLUw5iDdSkkXqRrSIHd/3ZfY12HpzpA/jgubEmaRIFUhOBJ2I19RaGN0qSTv5gd
sZl8AyU7Fi32kMv1IATX0s0w8keKCO7Z6cgc1Y6tP+LhNmUWpB2jHK2sy05rKoYL
ox0JoHFVn/OFvIC4mjL9fLslhIM+BjOKp0MfDDEEsj0KHkGfXb2ud+DkTD2n7DnD
VU6dH272N9KIHsE6jXMXbQ6485uw7d+1Aedf1iDGrDELzJ0yBVlmhjxkmBJBB63b
LUYKRxELSyPYhL9XmsVC+DxD/kCm5UFvWuIGaWLNXWAyIeACLVOG5DfZ7AEyz+N+
gUNxpWopyzxS9N4mH/iILTNEUNuEDVyfGXXjkaFY+nSTDeo/V9ON5MxaW0/Ce4YX
E/YY/kQrg+e7CzadDU/cwXcKq3ss//slTwzGE/EOzukH0+Tjyq5143PLFPNshOas
eedRUQU5nMEghv9Een/0dMYwpIiw+aqkJgFbIFpBlUI+emqtW4x2w1H149vb25M9
zSpkmzQry0WRKHVDv4ZBjD5drECiY/76YjPDso9oKC2HK2Tsl7gdPO5qDGf+5An+
pzL0+67kjZl8WJvB4I1zrpIEHnS0/GXhqdnma3QJCTIHaPazhHaHyvW7f+8yVLhZ
fMd4n+6ElcEt435jJM4IfGNvrDUtMpxDphR5/REZJXzhL5OYsyXy76drBDwkY+qM
TwfaviMDXftGWjfwPBdUqAkF+TpAiWnw0jyC07rXXMyOrMAULV+0SeemtEGoM5jc
3nyUf65pw2jjywMpRCWwXy7f/c+MYM3fDUeX6GCPQ7s5TL1LsCqKDtzxJXGTY9IZ
x4rvbvNySYEJqNSX3mc3o+xiM/lZm5IWj3CW9ZiQ4tgpbG3BNLcWwrsuCinQfaWY
BWQhdA82AqkQUHHP7O3suzAiPYbYzJs3NmU6dbp0F5Y4eaKnzTzV5/QSbKo0BIRf
87Ania2Au6mjk3hHirN4Q6EkR/QDUwORalFazUyMEPy9hCOLx2kgwS9QHfuLoEoo
jo2FxIywTfkE1zHHg++HMGBs0saHEXadWgg8BHh25Z5R1dwEjk2cQhwHU5KLKMlj
zhMJYScXdUEVvn0TBsgPUI+u8uUWy8fMGB7j59pIlhAMhh0F7d5qYzMHB6UtoL84
rChTEBTiR6a4yF6JLr5SK52lHBncNi3YqYGh9yXZShfbCaitsKOhfgbthrMrWcYP
Q3O21m+E63qiZux007r4WFN/0RKNYNrKBfESvvRWPgDqyGMwfnMbOrg/6TuDWWtE
DKKI11P1Uec/b/e1/7rOnPleV8ecEslv1NQZZNDeY+rrnOfma4GDac5TDrLASGra
gzLniXJYq/NYemVcjXWsj4HP9aDgRLWlMLjPddXgBkN9L9caJbQLKfEzpLGHPsGO
AVsDEp+/PtvSCMf99EKHkM+QCGRynggyxXa/Dz/cYmMHbsrQ82+LHxxjWHneJUVb
HdGWydsL5wegElIuhf62pt/cG8hivakjvP0ihIuLayMQ1MvMm518Ge+nsdZgVkn8
DBIG+TJX72MbLMMBfffDF+VUQzRsuqoEqn2+NJzhPgg30ITyBqLKq35hfHVDSgWx
oNDBP35PXh3Dsnh/UNnptX9WnCh4kXlJpFiC/FJdqGLEVgMh1yQrUfI9PAQ5oWFX
EQGCWQasBrB0x/xahgjMjjaxcq/9s1loPEdeRfZuxtfkwne6mVy1ighFy1d+Ovaq
VJUTqd2slaDp55sLlJfWoIf0vdQDCZNZisy2M9noodLYztTWqZiNwewfWtV1cQJx
9rgmxKvFeVRcv0GtyJcxQS0omSP+L8/r51E7oYbF0LDIpRxU0CZekuntKtoxP8e1
Cy2rq5BqpbXIVP35inK35FIl2+8Tb7MLV5tZmOl5GjnDl1K52t241q7FAj9ZyWcw
4kRRfpjyQX8cZxlED6/kseAo01RrRlr3bX9DL4b6kxMKtJ578jII8PnsKY2VAe2E
2A6DCh1DP9bs4NG74vTrk7/+Q25B6+tMBRHJcauT8ISVRIKFn3b01Oh/TR8RXC6m
6f7jFxkhF86Lz6kSgFVwuCEjJH13Q641eXmvm8Xrb48RDt1rCGDbkuORMZsFaqMo
e15yQIphSFPNs7l2gBx7VNqAZ9NqOBS7Sc+yKM7kjZhe/tgSAWAs9NF5F5537Gxi
aoinTBYKQ9zupjmF8KuYEDFJnQKW47U+yg718SBPmwiG+XvFYowF18z2yv3PzNT5
Rr/vDB97g6TSttMOUEmZBmttYXL3t9TGMRu8fHn1RitB6E8+R/DQqEbF1+OvPgF3
/2UT/05LE/tagUqNSzHcGsq69DaPFr8CwsqQsJgJGzbyjOlU51IYPsF45zDWIS/S
mHaCKZG0a4132T10xhwwMA3h/8tkELVdos6Vn8OCsatFbhdE4qVzJyED5nPVRhO2
R5vMzONdhjHcOjRh4euYibzZwI58mMGtR89BebKRtbWT2gr8mk0jAFtlHo1nO8eI
0wPfPOWBp+lkYjDag9bZsyq1D6p3gObjm7mRkOcn8ZTWi4xmfZCPmsv+B2oUiAPu
4LA/Q2jse4+opfX4TY7lQWFZRmDiBPkGd/WsnnwXk1IRcCK/SYVvwnVrDwtSoteG
21e19Jma7wtqz1TiB0q0cMy3TXzY4t6k71SVwtj1WUHqKrETwdZHgFhfBU6DJ0+Z
U2FU2DPhdvO2u4mC9D3w8AcpUyaWeoZGBVROG+tT9jfV5BTK2GomR4dPDJfo7n0l
7trbvXooAd4IQbE5jYPwUaf5Wn9nbC5jIyx9xTRZmXjgaSZqTROeHxPW9M6cj1F8
YaHuXfN69Awggx5hLBSUSpBiBLpC/Tfwn9562Kr+2DLS7uJCW3HD+2z3XqCYs1Lw
1jFGa16i/r7yiaDPusiETBFTqZI3JrPT0v56rbc886vNpaMAjq05iItXJM6aidJw
kh27J2wvAvm/XKsK95SFWobK20tTGelKOoBQLBw/5lrOcs3cIq5EXC7niXXQ37CF
lk4xZKXjzOg9aXP+vRcDFH2lnw7rSt/e3uhC43pO7hQ22Vxw2WRxAf/WqjMymUl9
LnJPRQqnL+zSZPAelyzjYaDi59Geu7BtWPjjxVd5O0ocYqNSceMQRhVJKJ2OQ2It
Ut1SLf0w+XbSsZC7CbDxiKvicQQbhvtSbJLKlWY2Q4KaEk+IPUPZxQbNC9PY3E+V
fKIcx6z9yLGrZqhJqmrEXu2IzlMKqsGNGzDJL+RyTQVxAj3lpN8Ead6dM+L2XVci
fOJVu7Q3hF7qQSa7DIUAHzkHFk3zvfE3Syw0C2xr9OOzQSS6WicVsnHU/F3z5d85
ye2sDjGYkQPrSj1ptQGmlxr4lNZiGjmZVtcxKL6rZTcb0Omx5qT8WzlKYzYCkRqc
/pWRc/hEuRaJd4ieqN5uE6UHiSPzo/w05H2DYF8j1ZFXULuKe2v/SA7Dgn6ycFKT
JmhLautonM0u9W2mrNEh0W1JaEeSTcvODRHDa79E8thgpg3ohsAb0eo93PfWLPnw
8ecum8QPdu20EnxS2nVzzSkZi7YF/KvSkBOS/yduX7nhaPF1Uu4AwMVDaPEdPWlb
Ykphox9aFDQLy1sxUNgUPLaOEIO7d4C1n1JH8c/4D0PaGn/CC4X4b322f872KNyv
b6GyAfejB8+9/k9kifiwhWCavPN57D9Z3W/RwWKO+tyTKL2MMT64uC3KkK5ERzxE
RzWhXLeF37EKGdn0U+pMMfzl+eBRJMc8xCgk7EBuj5tqjG4Vmt6b75gsocfQ8MTz
o+NcdB6pTe9wbsyubIbIhutnnh/LH1yVNhlpWQ8qHWaJdNmGjP3wIxCtdNh2ZMtH
ISDKIs1zTdVw0aTk9qDet+Z699zSju4frNu+A4ayrjt1bZj3tBcjW9snMo3czAak
rJl8voWbGe355Y56PEMyLvZJlalqr43mbaLIEveMzpKf5ux6SC+ohPhGuiqhquV9
YE+zv1B5QMybxryTgWZGp3rY0VrESMA+ZiZWS35I3baUIOj6V/wMrfltOttCIPNw
H8Lw9WO971A7DVjFBLYmEhDVduOxEwd544tIyFE/o0nuTIFCbEnqB1V7+/bdWk3R
8KsqQcjPPpNbCtRC8hhcUzvMVx7mja9pfqzmcXNLGoQ9alV8uxSY52YLihvxw5HO
/AGHklroSECXsXLFOhD2jTq9xZKowTTX/K8x+a5JHxVNTbgKBehOKfePQSqIMywE
rp1zKjzWxAv3RLqJz4RC1O72onRIwKVKxLeHJXCY8cHCWfeTRrwRhn+nKqCC7YgT
7g+61zdNamr2Dcs80yiC7XI9FjxMABA+DoGsVGOASzfUR5WsH6PUIUh0iUiMBqK5
6gRVHYooykGM8b+K/jgFjQX135WP6TsDvx744StSTEQn9Uwv7bwuvqaD+jlpH4A3
eTdJul1JI/f1npmBCT6T4ik8ATIAZyi9RVE5efVFRwAZ5LkOGbXJjko9YvUlA895
8xGjNyfR7L/kAeK/PLzKOqegwIH2dUBGuI9LLccfT5LITaUkquSX3stkj1oSIT62
t53lq5jPHH+FMiIC9FomldJ05fbBJtsIvf+7Oi5fkuQyB64A6W9ZAAhNc+ub7Q0N
NMqaCHPuEo+qRkjSr8a//FO3X51wGeKJHckz9aHSWn3CQRUd57X+R1TkThzK5KyW
sWIXavXbzmRotrfiO1Y7C4BODVpqZX5UMgyPpkzDP6bQn95VWZZ/ZT9BxvHCPHhQ
UxpfamMdo/giFu/S1rMCsoJ72a9VC7P63MzPBMGAq7TrUn2dMCOkIiZplMTWwYSb
g+bVyrd2DLD59IZ/Hr5LpngQ9a2dMGnNK5X3hOW4yrfOAHSDI1+GoAWtviKMCrS1
sAmh4Wgw9EvMW66+Ia5mTZFxCeTN3o2GP4FWoQulaBA/aYdX3s/aqf1w/RYaV3ai
fNQYOcnHASG3rPodR24n7BQi3VrVg2tgwdAUkCHbaUzqIcznH3z3Y0lvmEQ2Dveb
HaK4D5kRMFMVNtlhSNG+PM7CVrDTEAvpqbrk/+INWjtE88R1BQ+mG+yS1vu4DYFs
JuSFBm+BxPqFcS6vTFJVFDogajJ7x3ng2ZjPD3nbeJvOsYT4KWiIupNhP9mUiO/T
SnPvIRPtt8wjUcOIArBx0LEZcFrVretJCjSUNyCPNiXvI0P5JlG0qwu5zrXVDV9c
tZ3B6YQ+Mg6seo7HXzqMh5ER4ZaLoru35ErrgzYVfb9gAKomJ/E2U5gy/wiZQvKT
3UajjS3PSjcqxycBRwJrgAgYSUlP3pWMxc+ps2xRCxhV1f/4sTxGy9uAXZHPLWtz
JctLRAi1vdp/CZJsC81oAMTVeuqaw4REI1SYeTVLoWEIuQ7dvdCw1Cxx1zOKET1N
MRZ1LCflYxt3aHRYzq47t1w4Eb2a60+86+d3HBjCyu07PQ0YKNiSL0bRYfBoz6pm
Be88k0/kMvubgXt9IfkiG/8CTX99Ayl8WyUikQ1qX73b1S1ytWXJRf7dz78EnYL1
3FPWYuBNV9A4PFmKnGb/XH8lRDmBR+93jSs/nB+YS5b93VsuLRbdm+MFLJRmCMQj
AvTq0sIUnAriFrDbuZWbMQZ4V0YY+GT8UU3XZ/x3KgobCA0WW8vsfctK/FJNp93c
3zPCi1MAtC21CRofSWfMxjL7TMZIsWxSF/QtN2HCVU22wTVNYxz2oIaMyah6L1es
vWxKnV9RJfzLwSakCMS7fpLu8v5Q5Sbt8cYE8TjPM4wUrKB1r7nNiqQMMDhNC6X5
sKH4R0HiGbZzWQqZzloJLyPlv+5JwFWNLnDI/vqJkWep2JbsAbyPopNzI4q3nmO9
cYijggEkq+KC1jYq1tTEonii530KElqiGmL+J9HnwY42PzLY/34uD39C3Z2h2KcG
5czBg0zPpDZAQ3byTmsf6cANXqj5b4hkprTfKD0B2XAQVOPdwmokRu+ySA3TggU3
+Q87Fd33y54bq4BzXQsgIy4RYlQ5mij7c2oPHb1veMgy+vrkVtD0Wn1pw0JbZ87L
/v6v7/IlcO8sCDc5iFVjYfRWwVxqWzABanZ6tVRvHghFEyemonyMMRvhfLLAMMee
aYZGsMp579rBAKDve4k3aWAvXcp+BUvTgfd/iuy3GRHO1Ud2bqAM8T6VBxtRjyFM
6haLJy6UvyOSyMV2IL8/ByeInGsqVbPUrzj9Fa63JMvm7Fd0pBdO7Zax8KAtRsKZ
lvOJnWs3IlCTAF1YMFokDMtTkrw5i7Egda5RzAjL9FHzX7yK6awfa1bkaWxomspK
bMreUoT0oTPC1EXSYQ68utmNexYIDCwVQeS8wTZzwUn8C5BNsjyr53+7N3/MbDHZ
JddxvKuBJ6bRhgXUS/BtJWjVXaLXImuiO/C/Q1+rgwpvB6qaGknMfputOh9UNGuO
mE951/Eb+zMOVnkC/FV8WXlYpoAaEab2j9tDW38wQndYNt4+TPASp4RdnsVGCU3u
Q8W+jKmqI8ut+b6WM0Uv5C+ZPKk8wD7F2xwXoj2BiIhpaAHTb4viUfqy5mJY84Jc
0qNgTqPao390gT0PG0W6sMT7UYzAElz2mA+IJEyC0oAmQEJpk97HnXY/7ilUvstL
0+so1gAF7avNKfpkwmjr1whB1imQujUFh9h2NmSBXVBK3drJ9GzpEiNCyvFLQmEu
ZJ8ZCJNMFBWF4xJzku8eko3iWj9Xx4T0xl128kP+L4GWVYuEFXFMf7NKqQdAMMpA
mBC4qd3l8IiMr3gQt817jDtdSjrpmw+iJmQSDeghNh1K3x4UW8dNatFta9xpc/BZ
4EkZzrCQzoFLL+QZfV786rfurutqz9teUL1ZkWpKmKYvrPcHNY8jiLgv+AlK8kOE
u9TPmd5D9ZKaPf3k0PsCURCu+VOB+m4hGJ8ATZVZiHM1f99mGf6/B/5ELKTLbpu9
vZEL2WIoqOXtD9hXUIEL/NOQBrTKbLmDr1p1Zyc45/IrcOsNjQiVQGNlEoHNt4Pa
smWUJ34V8oJ3E0BzPcz8Rhw34d76PamL0mDN8MIKdnD0OzPAHMrkl+xsqUQTNlAb
huhBLkgrekbHRvbw+26LouRuciKgqpejWBbC+Lp7I/RkUFfVl/VPp6LqIqg0adfJ
oruAdrWRD9bj4AO8iGrmK/rWprAf09pmI6uB4o94A0rpqDwn0yA3PYrAgXGKmsIQ
4MICfQpuyKtTZZxBif8Ff3OKZ6IMs/sxVNninjDQl3jEQmBGesL/F5G9Zikt+8MZ
EeSrtqSZMLq7b1yEcuWdB0FsB/S/AhSBLe1zDO+uU3vWzDvAWENYOhNKgj9yRNRp
6Zy65PxXURKUuY6NCf1i8sKauN0mefWflJJNmUAfCpZViDJQL1LRT3uYPyAvG3YI
xHP6jrQ7kAEMTorK7MUFkNq+wiD/ORjC98yqya/8DmzBEriEDzc73AYpDNdESsMV
RhGw3jszhi2RqDw/fIQZSJPmFSJ44VpNQP3oDZovRPJXc7shSLr4ypt0JzF8uayI
9Tb27czpf483U2EKggAdrhF1tXi+jINRzTIsm//LQZiPH10NdrZsYdUVaQT+8pOf
GKKAO3DnvDmwtRPwsAN03o/Sy8veDFpIlOFk7S0UxexYRDRkwUj9AFIiAW829c04
ZytMM6GtsvL2POWNWvoB5/+mQfKd1jAMMjrzFrXcBR7NcC0ieEzvdecEgvHLeiss
RtmLLu1OZwJ1/3fpiRS7F4/1iBi+fJ48PQURG+TFlgMNarZKT+zgIa5whiOKbnW7
yaIbJH8jufQ7gP82yhvbJc7foVpv8u6JMLhfy1mSGbdY95eYiuLpQ2aeSvG01adG
jLGQ7PoX8/xEKVcnlxytXcZxmbPM3NIbUour572lGVbVUo1/C4WqRA0sQcNCflag
/LzKHD7GXGk9ji1mqSApGm1GZ3+ltCprMsGSmbMjrr4pbbV3Ww73Q1FS3Kgy7THV
qil4FI5GCqAamhifRa9wLXzrSEzIzUtzI0jO8J3J3oHpvexN/gpSbJemdcwt3l+g
rRrb+rPzmjQx4blHCoxGXZq+loy/XMPk42Q6Q+sE7JDMrESbdEKYIR/dcakQyy9g
3sl3H/T1RjF/kBMPmUAoX0BpIK5Pjajm07S/6MEFTjRO9WpWVN9khn8c/YUd+Su9
CLc8f3DPDq1hoc5eid9b/28QblBRWWxZQjB0npbbGrTZadHa59WIH57LT40Yu5VQ
aL12nhTuQRKWk2vYPBIcEP7AFhCSgVlCxQMsf8/Ll0A5g5ttmqb647QZih824oVV
V8g0RvvywXQkNi4sovhDv59gtnJDBE25qHOuydNAt3IdgrIajwGFxbcRfWHtgZUt
hn9949uXmOBOSee3faHugXLLiFW3o05wa9wmEXV8MscOB49jApQK+Dx+zzraFoa1
Qhf2zAZERYRHZ1a+Qe8aH9rp2ZrRgX/PUDUN6D7pEFB3xoJJYh3WhOf6MWoIellH
Zr7fb9NLg2VrsT3KgBfufLz/1/L/2nTruDJZgVX7dM9oUNX+0wDuGBlRWBQtwDk1
oF/HUgDKzys9EeB8aeyfnptJJd12UDF6jjYijofRbHeGDlZrM/YoJtmBuJVUt6W+
FfXom3JoSmFmqn4eKDJ6YiSnDh8qTi2mtdp57De08dNjwagwoUBNhE/H28VmoQ/L
FW6e2tNqcdshACRdVb1zpKerc9dOoD8DxFas3nLUucWPeei+N1lVGz5hB2vktvzO
e/T50PtgXI3/e2E6DKoM1LUoFGuYUz+4rE0Ozj2pVyMuKg2CCIveJjcfkFfXaOpl
s7NBtmmNSeyJkUJ8apsq/RSo6yvBw/c6UNOe5RSv56Qd/WhuKyf73FyuP2+Vldx5
Rz5t8ZCJphjIUYOEIUSfp1K+zCYpHZ+0CRrQphjN1rxCSk+VewpPknmqCS/WRHZO
ulKUKX/qafTOBtHxHsyD8ZFel6PFtg0g2dx9/B6z3RFuMi3fz4kdvypc9yKqsjUS
HCch5asWHv8io6Zag6xKlEJ0/aDl/1PrZhflT5P/BJxG/O7PRLHWp/1YbeX59/B4
wU9Zut9HdIMpbuHOf+g+E7qawk2WoMULBxwq5tg0M3m8L8kBhM4gT5C9hkH/oYRj
F0UxMEkR6iDd5z5bPZQSxrL86q7lvJ29048A0Oh+E6Sfj34HlazWgNP1u9HRS2rS
ord1iLAnnibcDZbAJQBtUw0bKShYaLhKwbywfx4KRY895aWv97Ar3T6U85yuJteZ
aaCWfRg14pbkYGFfZ1rv+N+j+irfR5fLmmEJBpM3TT0/uNSifn/UDnPKFOXdl1fW
DpMxs44Rw2wKckL3lBUlfVoDzOj9nOlwfDslZVZiNQyFw4PojvG2LNK7IJPAKpRd
mbme9aAaDMT78RzGqOWhbKfEaMge4r4CktjG60jj3H9ovUhqxq2b3cDe5bkCDwm7
egUTykVWTdr0HDHOhL0BqVrn4OKVvqQJhwKqs7YN9PsLnET3qNeLsUcSRotuu9GV
mz+NsOU4Gl29bb04nmJOr3IlPbP8bS2pQM7v0UBil6PMJ8spVsM20GsVARtArF7f
fqOazaAlYEcMTMDffeRpvx6Kr+kF/qRta1QfZQ9KJ/j4epN3z2IZpPRi6Y9+4kpb
f7nQHoaZD+LKSK7sTw2u/WToeNjNS6/sC7hUFMJI1MZobdloAeud0ylTtib4pUWi
ayWF/RwhrKBZ+SDkFMsuu5PMS9YgznsgGQnGmJe8QmywCXw3nw6LGj6JV/zUs3B2
VdXPum6jjsKQmPmojkl/aObTAGJTq3FvkHkv5iuimmo7V9OrSRjePazbwE/Q3qQs
6KYkJOzcysDMcN60gnOedybAYxxXZMswB4FJPLVP0fSlMcW2OPDQsZUjgafBn3d/
TgqBiGwW0avKtAoyFLRG2qwFHxnAPXQmZVt5nqgmCaKTowQjIyWq7qZdnvWGW83M
VYDzOFuQfW+5JzKClP5M7xclUto6eNBOHMwlyujwFfmO+YHMWNpHk1LV3Cwoso4A
+bwKWtqBCgfvtH7xVpcu+WkT+SWvf0fl1s789lwmQm1bAB/F3sXiC8PcyMgZCIK/
L8bVmzezQYVXQOAip/nQ107i9VuAne8xqgaVn16/9cTO2Sfsaaw1IyoNEq+gHaFN
95A4BZR3WgyLOfUvED688vFzeqPxkW9P3v6tep+1WasU0gSyLoqxtuiODDGMid8f
/3IkUkP6X4keCAXaFVZ4QVpJiwN3rVZJbTwg907fKwQvskIzjm93ibe3w6Lk8mm2
mPOD5zZeprJbTkIEIScE+XW1baj5xXXQ2x13ubG9B25f80PmJUHBAWITU8igDyzV
cglW6iyvvZR7hFRNqEpQwCz8P16vy4kLbyxiIkeHALISEKQEGSK9prVh1/lHOsr0
RROrWj/6vc7MlEg7PUKrtxW+T0GEBQlv2ocl/bq+QFl3xDK8a+GYuYw3nss9eJwh
WhaeIWvU9X+WXFpxAgo2g+NWPqNH5jnPou8EZnQvuQ9IG9iefo3MYyHoybAngbdy
gSsK4EKPhEQUL+t2h5gMu00+A8dJnXgDaZRqk3nYmZ59GHsK7cQR3qkeM6Lwom4+
z/xCPwhVxnY2LJdrwAvNNRcKS6DCkhrM4tVMIsJsS8GAeRYLt1atb5ZZCrML0mRK
imTL/B4EyARyuMbicECGh3q0H94NGuEHWiskzlE4vRvUAelolzwIIdj7hIwb9jBl
pQPjmu5xfBAElBOTntcNNfGp2kQ2v+FKGPV2a0sZNe+XGGNRUxw4vutd7DsRQPvW
gScaV/9E9khzxeeKQ2eEMgvbSrvxtwBvyoIQNweGWV6pfyBf8Z8hm+tNEIS2KaHa
ogo5ArAq8P1TSVcw6QbqNgZdtYPFRXeUONWuEAyHstFyzffx7213DIUtmqtABh1S
tIUvCUW+BwN/R1/UjqV8IPay1t85zZ25AGvjrcOrIXOVpxxysklBDIH7cuc56SyT
V1kZo8OI2Mr13ZIUj2QFMeSHV0V3aLzSt9CdF42RYklRaf2iA7NlxP3n55mBFRht
9rTPtpMHYxNRWYKIIJec7+7Z7zH96sC4gsNfwFO8SsJTzD8sfdHERd6lPe7pflY3
gJX8bCb5NTM5T9wQkK3D6iGP2GTUYLQ2IY5Xjtek0medFCQJiu6gXzdhsvzI6687
Ppe1G3LErl2oPSuogZwbgSjlos2NpNessJ2kPYCnmr+5cK8iFsitv+g5OwkmLWzq
V/nugEll/4nSEee9yjMc/nRnEiBUIw2ECNXaM1oYi0dEtn5iOznfkrasExsM/X+h
n5WiV67P4GhxE51axL/3aue9gZm/v+MamafRyaQx0dU0htTBZCleBal4zSavwAun
fC/BYPdTi/KI++qtofo1oqVCC9JK6nQjuVaYEW/bKijHBhbgCoPlzl4lo34OzoAL
Hbst9gNpoUzyzlm0RgjuP0CBR6Fe0OL81aMFlAVEnfJdlP6gS3Z2Q3La9j96gAU4
vLe0D7QsGDx2LLObGLONThh5e3dLgtw/YjqVZwW9DKM6NxXGTh3QazM/fyfpF/PC
pce8QqkhKA09COmpAm8Ok0vAv/tLkyIt7+T0WvcR9SsYjY7gzZr2MXiuTYUWkn3e
nXnyToFjkhoOZNCScuWFSHNVu8tv3al6aKrjjmP2BZHFkZAmT13wcGqII8byuJ+I
BZ2lhbSGzq3zU4+9bnWnCv+eWo8aw+Torxf6MsGgJ8QqFGN/sdJSVcM3AdVs4ijv
zJfQNbOm+GMzwWA5PfrRPEDwl2J326r6sBwVLvNAlh74SWJEwQ7iOBk8/NztHTqi
/6KVap1CV+QIvImclZ6w9FL0Fw4n5oUgBuYqTGLL7f4RTdMxloGef2Uyk3OdT4hN
n84Cem37nYj4hfXd7asmLS5mY4s12/T3pQjRB/DyW48XfpPIMPdZaedvzC2MV4r3
xac1Pqsdc4SQH6AxrSD5RCRXB8Cq1CjAU9VYn97JDtSTQwnGyAwRXSoESj1jGmkb
8hOar0B/RCm6bXIClard74Nj2E17zf1fi5Yoe3AdM+N+ej2z1s5preajTVW+02RR
mTY/nJowpd/cE7EYDaARefC5CP3CrKGULnRjzbvctlGYiWsMSbgynMcNzaW6hTvJ
RjEv78ltPDsv4AUzY9HDiT/9ziVNWv6XEHTzpAwdjOjWv3xkca0ziNVx0zWF3iGD
2ura4xIlknFFR8nBFRoTq751mtsSfr0/WDc4wwQUBpZRnr9pVw6WOqUwYYGBR2sd
eywSGULpfVaGRQojPacmzgWozLMysfpAZNz1R8vChF7EV8HQNVts8HZBbsqkGbod
2EoCKKV9De7jxkmcDbzbaVTFynfVJ7VaMCHoIOSTb9iZ3hgdu+ZwE5qgL8m5sejp
kqXN4IpYRHJf1Q+M83AbnMR6Wv3D9nubosiUWDgBeFAmhJjOujPwv6TnIOif+xQw
pm1pLnVpIXqTK5tB7j9O9cOU4NvHwenla2vFd79JHwniE2R1BrfRNXqZPkVY8cAD
WsU3FJ4jLAaEgPvlsu9Oe6Fk+sF/bFd6D6AQJFHPC39/aqgGNR1bW9JKSEvYgCGm
dpEtBYw2PnUnkt6MIlEYgMu6z6lnsP5EEi3uelF2VXANpngK18rC21FbXqhdg9AP
lTb8r+hO40C3/N19izbHbbYcakFoYFLLwSUF0dadSKfG8CXVSd34LDlfhpk2ZxEc
MbL7RPiKaVCt7Ejtz0k76fsvWIkvMVB1rT3noTgM+/gxXUdPm2RUcTsVfgxjgTws
OVwjN1FPahMlEZCalE8BlYdeivDnLXBxJF7eMs6HFhoeHSZxxhr5t3tbZOtZ3K89
TQqUNR0tJvrcuBr0R6bHtt+I6TCw9Je/oV+DBudU425x8rgAOHCgS73auq2FV8rT
PvaWIvSEJn8+L/mIqHgVqy8LUfMIHuHrjel4FaAQ6ym6x7OmL8/evptN4YoPLuGF
yTUHAG8+tl2UkKIJr+WGPgY800VXv64v39UNUXpMfdfNo7Py2uW8NPy9D/9axmGJ
z+VX7zo0sjm9KLLSRCn7MC6a7+MpaN3Re5BYaA8LvfwUANURGueAODb5iEgxLvQt
DbgXhuOEJ0FsixfmlWAQLcxfhfKxv0rA+ZGG+qAEahLVsubOFgzhdTF5Ub/kNRR9
hHnEZyGR29Fvyw4oX/l8to5Pt5S7hxwZ8IFwM4zDYvj7y1dg+0HCqdhMREctzYAz
z2+SSp1q0l8OEq5HEf2Ad2xzGkfxL9VgKXAQaJ11XYhNWl8QC6+pQ30pmwo5rtl/
5FOWq07ppt5cyis8rLbNdYKDGh80Zm8dHCCVfkMS7waFqk6CkxorUfeqaFP1rZ3T
USPN7pOo93woj6k/f8KxziKNdF3lHXeXWKr7SrtMoeyk2uBChINKb+sRoLmZrKQ2
konrRhgdQf4zqu8LRhVKv0VUOGZXvX5dDNlsk67O6SBc9taTo2hXLxTlRsChVS8D
xobul9GWEClrUZi+lSLWzIjuD0H0Oz2TXbwKCv9FRlmAUz9lNJLoIfv8g9hw6YpQ
lRxCbODXzNXcQGbvXz3K6CW/FeWBCp88o2zmwGseE/wFc1Dv24en4KjSnH8m4uCw
J/nND3L95xPNs5EF8QvfcOK48FJ4XRJkD1/yAhH6mTE=
`protect end_protected
