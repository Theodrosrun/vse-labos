`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
WyiDWudFU3KQZaZWl/rKQwSvwPOgp/YSPeLOMGuubHlsT7JtUCEw7kONy51uTO3w
klVHDjyZqj/CT1R8a5GLdPQbjrhsIhXYuBQYA1aTULzxZppxQmOfpbMekum9TgrO
izcMXMRT9yVx/95fBa6dySMOJrHjvGZfIKhRhTql8e2uPGml85tN3f32DYDZyNbU
WLPVgIdunWxXggKuOvvdEmJkEzwhuzHaRBHFQJOMxGLFZFgP8emzEPcC1EX4/mEP
uY9wqphR+zx9VlpVvIKxCm3BjbZ0BygnIwiNto45fk+nPTh7AKORXn8aCtbPA+AL
+y8qpMud9oah80FGyPhtuw==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11232 )
`protect data_block
T0gB1A/4c/lw5wA9rXzhnlBJ/ryHCV/jjS34nRHei7x8o8JUbCBaoTd1hNFnOuPt
MttTjf4lrwzEkI5SkJa54hQLhhUYyPAZcgoku54nEeom8qqUnhDvRgFlqemlb3eQ
Maa3OPngAwFBEV10jhzNm2sfP76CScGZlVo8jax2h/Sub/UjYFntsUvVjvghpqHY
qL4Cl4+tkrn+stGBXg+LXnjtkuGm3kNIRsm0NKCIQFc82yf6egWYEu+B3H+Aaeun
k8e44iN4ESffPdsDG036YBOI00e55SPGMa5+sZCzkou+9P10MZ76ULIuZiy3rOxG
9L9Ktevdj4sL45aMp2jl3dobRQ2W3pKIIzciB1/kjXzrauvpk4dv6qUsteCZPP1s
0zlE0TVgPsw+Hom/8CJaOCr5RwcSPE4KOH2PX1cln0gMQs+DEkbl2KbxIkC5PcdD
XJPMhX8e/tYunaGNzsmZyBkNpbGLV64MNRlgK7rOk7KFav1ID8sAfPBl9L66Oo88
Fj+c76SGytwPqeHCeyjS342qGTDBePQgfaJI6XZV9zK6QdFjjbQAqvLFDLySznyr
6vd6mboqfe5R95gu0Xhppvs4p0qU/QHvuV2o14L3POAjDcxKMQJ6ZkC12JaJKhEZ
UlkCbtoiYbENGWgls1SVjm6WdKwJRrlXch5lg2A1vL9zBKpKiT6f+l8eC4XmvQMC
XU2xQntT98rsqGn+TSURrTQ5MLd1DSJ/UH2XgI5+KJV7iFcTmyI32yC1COrIGZHI
XNZHOLAF+jh+q+27B1Jq1IEzCXw51sbwGJh4kYZwnicqyKJsgcqBMP9ceKJr856X
9lqvpfILVucogkAOAKS3nRvV9QLNg2xacDDF8f2gRf6+Qp5OJvl2sTR/2DnzpvKP
XTRvoGNtTVoqeFefSc2NJrfxEudOx/AtfPUC4H8sK6Jvyl2JGac0pZ3XFHmv5RYN
STuAT7M+V/BAtGD4Bff54ZXHY90VCoyCnwuK3V8UPp1JxkJwwvsRTQtvld9CRzuV
qNcxzxWeJhGdCLLpoqDi8UmnhIGopXPCfbuQWnZ6KVhkn8b2mdSZo18MwjHH1Ldr
Ahpk3DWW7Lf7+28J2eGH2fPzLd7CYawRBLSmMgvX3fHz3Avi3Bx1scYTSpZdwMl2
TrmW8dbx4czs0/k5oIIM9q3MwBEORnXh/6cQzQ44XTGua0VHHsOSDvlgWcRXHmZd
G7Irj4DDq2vnQ9nnqU69/K/vG6LTgrT9t6oinmQ5rIsd0efBPyHTfNeb+IRNWygJ
tdtZAQzyrI5ivS0Ljhi5wunRdxeQzbAa078Qjj887pNB7M0W0WZ+KZI10I4dBYZI
tLuMURhWQHCtRWzQCnYNX6wHe8rRsjns8XjXVZun8Jmr2f5Kai4u3Z9noI9onK95
hbAvJapVCCU+rpsJXCrqJK5/J7RULUMzzZUMGJIQS8TBQwS1/4PWqAzMqh7wf/Po
EJTrrbv0EkJwdP/TQFVWyFtr9gnowhsbI4o6S86oqrB9D23FGHRMgpm4ZRvlde54
s8QBPZd03dHyaP8D2MALNuvjLQUG82rqkkIbkteh2XsSYI3yaEX8U+oCnNyaoD3d
41L7Q+82hm9OdkWymgAL+sWjhsSyumd+YNBNhHxZtCfNlXxeSd6cpoc+81SvctRI
hu2o2ZTEA8b9Dnnxm5+QwAmCB0OLb+1LQ5zMNjSrglDr+l4SOURG485tvijEonkA
b7nlbjYsDC817v9/ojALWcU3WEMKw1V/L56fEVwpJbWMnNhnAAS4dysVmtHMYZAc
t9UwRh38QGApdG4G6bmx1f0EwtG4vl+ZzwFtPm4F2fw527wZMzTXsSBhrunBmf3H
88V1njTTM/76bpQ9/EnocXXkmqlg12siQqOKjZqgp8VO2KbhhgHSj97oydMIFBC3
mC74Eb1TiUneLthbkJlZ+d6Hcd+g+H/Wh19RQ73T7qeBGPDLOqnTZ4D49SUhFY0Z
0DWOwUbIQmlZHL2CNu+aj4PtClYVJ48BScL+Af2p1BkkQVmXYZH+q/zDIc1K5Oe8
4qlnS2OAyv5Q5RAS++HgP2imAW6KF5wPFZmEFeS/2kKlEzzSse8rWy6gxscunf6R
d1gudJJRAyKuj1ugomUC/CPjy3f5OESHvFyrBaVQ9XNpmhXqDRnbdY2CHCrPs5ae
0X2p6H+rffgK3Jh2BB8+XbzybkMt6j7OKHaHopdWtv+j6/CHxKtoxkw1kq1UVSTA
63qiQgYWZ5j5Vrq+VM2rDh1rGrn3sunfZcGQVoDZ3r5kY3EcVRLXp9/0qBYcVwI7
G5eW9DGIOIS2K/2r5Sv3+WJr11uwbvR5ZavIfPwcsaHnBuNWzgFbUn6TY5RFdf/J
HN8joP4ID7fsH12Ug5wIcCHSJbNo3vuVvtGkIIvibkWIIkOGkvZgxITsCIJ9/XWv
qXQnk/jPhufVt3neBw/dr5r193XTxuGv1tR+dLkFUujtvjczLWU56AZUUiNtsig5
oTeKFf27vJ4KQ/zcr4nAeCJlwxd5hLlBoX9tzpJza6bhovyOAB94dHvNS09PaHyl
UNRiuJ0CJgGFo4VuFgL6JrNE7Nb8Bg4NyO29Sxyj/hSb3yNpHe2NmijY7gl7Pw4j
NGPc3M7Jy1MTGKR7ylBqPBBed3vNv5gttFQKUOMFZ9MZxtRx3o3e4ii21tQUm+AV
Est3kXXnO1N9oK+OEtc9NtW8LuhsELNByGyS2ULVM/W8N2rdHWkW32+z0qmTv2Bl
FlZBaYFbwZQwEGNHmtAOgHAqsCy7oOxCPEeUa/49T/1cbiBhPPF2XSdNJAwCbiiv
jqdAHQz8YrHzIaW8sj8j5q2BCMNR5pFqeT3Y8t7v5k5eqT8eerscvURUMbK4SXDo
1ytERruDwgnaV3x8FilqwU4Vs0tZw5CAKs0DiO5asG5nEiNQ0wEeO+gUDfRj3btu
5FGWgMB74MBfozaA5dKq9785iJxM9Mzxwpb0Q08NAyTsOHblqiXbLl4/599S66yf
u7IceUHfb1dCUSpu4oiAmZtTYVHVaR6z8xq7CKO+YRARyqz8nDpmdLVLPPWaXRlg
ET4HthTCBQcxtrtGfydldY6r45BGSVyJjL6Kw/afHjIUomvFSreGggaRQ3q+QVtX
5njdLmM2nQBff3vWGKlW6IccIU5vgk1DKShji7ZkgQawYH6+8WwgEowCWn6FOVVA
PPRTkYBz380NeN5jvpUzsWk6ePqnBin4/eePBkvhlIb33UWFNXcGjBKSevVRBDzK
oWHe+mwHsdR5urmpfNazRdZW1z80YwkDk1IvXaHhLfMdVPbAn240lkUs4O3VdsLd
KSnEZaBSWmhru+tOGHtAVUg6hlzM4eRSbl/jWri4jKtf0RM6mT93enzJHno8PRst
Ks5ehPYqgs+rh0uo8hVFA16Nn+kxUTUKSU04gRcrs9VhJeFkmJyATqLAzhvRmSMK
31+3BDp1oSnW77sYU/L0EghnbP9eWtWdkx32IXddzGUYbAFSU9X/0OQdUUKY2P4r
bpDK9mKykbcy8KxHzS9wDtTbdZ3VYaNkXUFMFlF1Wo4P3DN7Ycg4b8QxkoNsGNHl
PnBu8a0uaJCm8hn3lgfCJl4exJHF0h1IUYPyh7tjoOT4Ji8LPRVdonZ5xSGml5rL
uzfYY13IB6rz2ODFurlCpmfG2JGRAgUQJQzdNjgjyT+0gWE+KA4C2EuxwHuWIJAA
vHPWUfuHcqc8b5p98kXRRcPYeAWdDHBQ5GnmbveVQLYouLCZS11LNGlrmt8r9djg
fVrvwX41tiDBuAxuFPVF3fOnBHs1rMn6euk+Ssl4L9514lXAxpL+qB873rC2euU2
Ivo0+NheTHB1lpdfhuaXLM5AHk9FMW6/pdnpF6gPmrJ/84z7H+80b9bRHsAA7nyl
4TbZ8OoCNQs2r3HwjR0yek+A3pYcAHi9BX1AQe3kSTGeXMD2vF9DRGXavtrFLWeh
PmMu4GU8n6qswLrw85KEH3kce5HyZnl//JRYoI/JdMqpmPeeN8IRSNg7LUuY9/SE
BtlqN3YhWlxgGOvka7ET+IbVGOXCYG8uk1BF6LpFYmfOylip7Y/jY85x/gWV+1JG
5hCtCA67eHhAMV/zLypPOAgK4NSNMIo1g7mQFzrZo5S425c0Qv6JtNwZlAXBfkte
y0V8D5cnUNrn5o2kCMjpiXA1vunKGs3h+j3OW0019GNtTKvlE2NlLV802tmyBNVb
Uinn2OYSkXpiEaVuspfuNzclo4ICBfK3iNJVe1+3ezkUeRSKCfRkIPYBaRAu+FtN
xNJcvnl7M32Nqm8muiOCNuEG5nXi2HgZekqlVhBEeHejmZQt+O40ASnpUrO8MyGU
6ad/GPht6Hyc2l13Ui2tlGzmV+hIZWc8GAIVTjkd6p0Q6wK3VqoXgjrCpcF4ds3L
q1jKO7DPIh/8YNDZQ01l3cyKwPPxIMqKqpomMf5vzkgLOFq15KmBAD143k78vp3J
P622qa7ARfunFUb9jZGyBPlI0XGqM6sO8iHlExh2HS3wHriv92Xw4WVn6ptVHNou
voRIDxbEi5ZwR6nFcH/UwUBi9OY5TBOwEGr6teC9x73U4frUcFlDagZZlwvxfAZc
7fFjMNV4mKk7WmTbOvEhFyWiokWWfSC05qwpTdIl0sYQyXRrfZudZXcAZpXG9OrF
cFmdovH7jhHooKLwYQhgMRLCUaTt0kDMLNcj8syPrri3sU5YJd+2ZVrDccSpIOiA
j/1OsE+wxR0Y6i40dVMAmP3d8on+4xYS6bTnfkR8yqEdlCPVSYNfccgCFZs7SMhP
tsvRx8G3KsfZXL6wN6bE/+XSvL1lnIizf0493gAgQik5A8t3dvrx6surYX22Cxsu
GaJYy4fPC9rP8ghoU5GnyW1yj6leVb603lYGWwcM1H+Jc3ht5gZlTtwyxID045MN
qc2/hvR8FwjAi84OzsJXAf8I32F7YoJV601PxRVz/YMNHsn0KzzeKMioAeC1F9Ge
hWoYtqb5/RboXg5mPS36gw7mDVZZSM0uGFJD8MMqCHStEbms2OvXM3B6UVywO2SJ
mwQS89EYJkiLnN/5jh30wy9cWM3dhbN7IPPpF9RL6YQTpwAED1bDdSSMWv74Ase4
R4eNmNShRoxj4OxdEJn3AZwt+426O7+89yiQpItTNJ3rjSKBS/17UcX5Xw+cKBkm
31dzh5yoq1lcEMhgKp8bUSn771C7qOvSAg4u3f9tGQEajrfilpr/99TNOeI+1Ic1
L5Kc49fmsrH535ceQO3H0C+18STZGJFlxBRQM20bZdMFgBry97K5FRfx6mC3FhQY
OYoPSFE762tX6XI0mYhLfOLh1mVAQ6zh92TAZCK6pEwArAQ4Yakdi6viqCr+dBQT
3qN8tUDYMAVvX4H/LOJTpS5VtL38N5MF+v/UtVzzYhBswQz8xfZyWklkz+Osc/wI
GgEtC9DZxdg5LdPqFrpWEVha2pgnhrZPIjaAqAjf8lUpjlTJWpyYwBZGi7b0MWJ7
vUNO7CSoyluFy4Dl7QyDsFBs4fmtd6lEmtSqvYD9VtACdnbbOTmN+c+F7gucyBK1
Ilv7PinYjmtwGhLf6P7ETmaOR8MWuv+egXDMv3pg4Ho9MhLx9RARydKqKPN2Dzng
AiWCnmLWGUbLNjR8LYSPZctS104fSCQLdxEy44Zq/0KM+D/ZVQxSfF6UCtJlVwKA
mdahJhTEZ+/ArE6EszfDSctCJC+/kzZ25fGUqfuhln9PnzBOAPpkUEhpERPkZKb4
nuUUMTPDMy4pDwuELDAxuQ//PzXkNdA3+zvZQMxlr91NTiMNEA1Rx4rvRKG9jb8A
E8stY/hB/ZTEDYuGCA955oCoPJWNp0XPbyRht1Cq8IzDMra/1Q7kUHecA44cdZNS
FG9MtmmbyaKPg3f4TzYi+QpkOkiAyY6RbYy+GRsYqcoiP385gTmz0iL0sFZjVGYe
CHC3KtHn2/PvJgFgTmAV5wrT5ctUIkE60UPPQLtA4d5dEpicIYB9oN6wwaT+00H+
07vL79Gh4c2oK9lVrrvGgdbDa0sREoJYLMItlz5Ppi1yu1CvZpn+o3u222Xp1Bnv
SXxfN+dd9lM6vmoCu9SuHbxjbe41EljznZ4CoEAV6UU4MBeVtmjKaRF4c4vuyJAa
16sSYwNc0LDsw8jcjTBu9DvDoYwvX6JfTxNXB3vkQyucn45rc1Zx/RUYdwoPJa+3
V6PqSq7RuBO9pnLr0mrqAj8lc416cXI2wm2g9krLm8KGqJWi9D2Vr2pxg6zO0jyq
tzXzqPrAAPJPcRsb0ZtKQldIWxmHLXlSSHHbI25p9Mk6KwP2iSWrNmYjvMDylqTt
LJ4Kx6+1gsmdPICcSLq+XS63PcKWB1y7GK9YpeEbZgtkCQBmWJnrXwTLzgZItxYx
JHo2qB6KzAHACwczabVww2jzS6XuhBsUIILVxk9BxM/0bkqexx/KcFiXPl1UlDN4
W7Q8KmzdBXjf2iYP68/o11k6tb2uYzCNSQ8U4lQkJeal3gEnIuMer7OAEQJUHhTP
TegBkC0JmGKFQBY5afLEYXjSRevtgH+CRw75sy4XDShD28gBQ7XY1CFXEubSoVNe
I/4Qlre0/Ina01SxS2WLkf+53aJKKtKp5kftlyl4yUVmwnlxuBNCwR04QubIdOJ3
Vg8uxH4qpq6DSM+NHsAOBIUqdU+Vwuo7Qp49xOSZ6bTd/UhESZdvSQ3ItqBE5FKP
QaJEeJhshSoTp2BFQJQ8XXu24abbgOdqsa95Bpm4Z+hJ7x1Csl8/QDDxFVswgqad
LOVukqdJ7v+znZnM5ItUnFVM4VRQajsOiHcK0FIh31/1WOcNLrGerGqfWdZRDOWI
mmyj2u8lFwORAbxkpVVWpMKbWijKAQN3P+OHDnRle3+XcgcZ66Rzt/s41UVv21j/
fZy9t9LwP4fqkXvlSn4Y3szbIWILdniq+qEkjawy1FXf2t/xrRp+mE2rKDEqN/DA
OiUwL05c5nzYmKt+LdVhseU18aByedXlcrHzrkUqjFr40dAae7SQ8HnswQ2bDFaZ
FEwr4CRJVJxUBLpJ07MiC6gXNz6pc2DaQfiw8zNzyJq+nFWbYnxovLRyUJ5dbMdL
DnankvzPyPnEZdW7IG7Ul7vX6SPFjKHCJB+0H6h8yFRyst54ejLfKX6AJsRsFKBr
GUTCAx+6DmxQWX994uIGRzSmDHT3CEAL4/kMGnVbmd8fkSpf3JK/ylC+gY4puevZ
DZ4VepDh2hwDojzLTnGP5tpNBSkS+NSQGz0/2+EipM6o4P/nSYREpDH3D85ez/2y
xQoqXpTs26sD3FyUpOR015xdZ9qtYANVZ87Z+S40IwUtKodg6E+yajsO1FeAINAS
crilTtwaP/FYz4jn6MGEe7ERl46rFU/zio97CTkuyfuQFsHj2aIg8rP8nCfQpNRk
cY2RduWEXOmuKnI/LqZF3RvjHY1A+u90WiXt5qpmcBgRYvjKpKt5RWoZnu0pQu6Q
MrAsBVmSjhD9LKQ2uA6m5Ry4OWzm0KLS64FDn4Y9ABqejtzpDsKyIduDIxnfCm3I
g1Z3stmzwhnh+JXqq2yiBS8Ra0+Y2XkUmnTMyYBpGzeRvxx7QAX4UOcQxzqi6wUE
7QFeXMC5EAHSNRTpr7D4GIu28Qpo1pAsQRyloaOvBSKRmZcs1b5Niypf+bB+b/X8
e2RcjaLUqFqkPaUtk6gMv1U0NroDmLrtrWi5gEKK5OpIVmT7VltzkuE0aZ+I/3Tq
GvU6nbMbtfIqUl9M1fz34VvGbZjdAnr/CbKVgofdRFFsHjfWMJrdNOUIsGIQhy2Q
ACW65dpGBaCmx6No8B3IjMpSEI2CqO0hOxyv88nZ2M0c/jSXwX3USglvkw9LQfUC
cwO//c6qVPHbOYNgAooVzkqo6WX6IODKExr2TkVUMU+XDiZ7C7qLKBzKQDPKPK6h
HxxEcja6EgLR51a7l2iYp+LnrhIQxaMcYXYtNL4REhiXwlARHu9QpiuKg388gCAN
qL3UAm45iyQgkgoyEbpNdRqwZE3pjjQaZvzzyW1IbjL/EdV+6VZs7W8d4BbypsHp
q0vCLr71njI6dfv0GcCBeAstvtbTpKghEE7B9hM8x5lf0rFUvapnANNcINkOwX3Y
Kydf3gIkvIHXgHIgntDDIXyPSn9golaUMeNsmOqch8mi5X7tHFexMmHEGb9gSp2l
ALY6//fNHTJZkdlb/PsNizXN2EQZPl2IrsERsO3+ys9hbbtW/Hqivj0lfVjvwoGz
ONJ4NXXmCLh8HkD/FL6a2NExuTWyBiQK5iFT+SvXmwaN1CVhPXHxxW1AlBzShqOV
PXvTyPGPRQRCGSkS/4Mk5FIj6FLFex8k4CNFmYdCoETwT8DnpqUqAENuUMiYQoen
IqT0g50H0EwSL8i646JMRP23GMyIs4fDuGFgKfp5hzPVNUu8GQvadYZjVcuBUSsx
t1Pr6fDfss+qmG26K03hUSCErrgOCUZ3E3kdy6NlkFsPm++pDhsyhAHYSTtKCONv
R5vgjrB0YhjgBg849ZIAmotXK50D9iGIand8PmfyBUCNwu41yYF7C0F5R+H9ksC9
v+cylDNhiJVd6EZjN4W6wwMLlgSH1hwPyOr4u01K0RFepwaZS75BgJRFXlFmebkO
3sHjRroZ6R3YZBynLH+zkCyc5OLyN7eyX5+K4Aey3B2zZNSOPQXYOEHQoKlby0Hr
4ifLeZapUkfAJ9fDQf6Ki+KgmR1McDwrDNA/YnxwJX9QTE605TqiWS4VsdGit/Hg
w8GmGeSfP1ILV+1HxM8J1SiM+C9EWfE+zRpI96FWhEKa+0uBGLKDs6lGkyxAkSsI
9W1ICF+t/PJZbcQCZBl9/Sy9DRROKSEfG9SFJztIhRlfoTbVmfC0OEQagL6Vn+Aw
0/Ixm3UCj92hlQJispr++6C4YuwhyIGASEedRPFadbEIUIO3G8cVPxFsgVcsP0Gi
1j98585/nkUddc8NFyy2dKqSnsKXrBWD/nYeQ1fmm8MbksMV/5sKK0a3ZhJLcnr/
4r/vf2OLSjcRyiI8y1yEC8lvLtgaO5N/JQSMykEGDnZv+nYTDvK0Iz8lZA4pVwlL
vd+KEYePjdNoofBx0jEpcxIMCNkm0nRr6vd6ZjctdFsXmtw5rqk0l6tthkccLoCc
GzG2a+reYZMcLwQmJm4sdbY7zMrecDLxvtK/ixepmLFXdEYjl/TIZhjaZX8LTFq+
YM6NM6ho0Lxe/uCbjXig5pacoQFh+1NgPDDbybmkicSdXPu8WlLWG7J5zdEUWpc4
j5i1h2wrPiEOLLhtujK1AVgVupsjurMZEtGKq92oi4h2POx/jVFZMUxlZUPCuFcg
JYA3E7H+jObZvjW/ogN3Sn3kJ1lPBmGOib5n8cAWro9fxEZvk2i6/I4HCQx9U6kq
eGIr0KCHQk751ZFkUB3FpHIXualFQrnf4rMxxZKiY1A49gY/keDDWgC1EEeliNwC
WbOhK4PvreagfgfKqziJLEMtnshYgyYvmWZopW5XOzgcz99FJRb5jcSApqVn4I+0
VLU4TNb3+HxGoE1TewE6vpuLUViwqZCsR6r4Y+5Nuzj9wEhYF56eGfw7Dt0EAXiW
Krv5pZE2CdlEk1ip8XD2v2kZXbbrQYfd4Z7hnewZdt3HrEIHRlDMKf0rNg52u/+a
0O4I2QZyLu3Caq4d4mCtHN+UCwE3XJ3ayohu4Dzt4PFGRfm/0hE/gKnyLeJKICtP
Mdsytc2cUkhzFluaeblyQ5A4snUgMyPciNcHlTpoEbxJlhmRuJYGH+kzcyMDt8BL
1sUjAy6/+0FYbkeKjetAKGNS99XJSzm/OBJpL14h9AZ7G+SUdfmdbygmnN2vL5y5
5iJD4xdjjrvYpxczjOii2qwY+7mAe9wVVLK9A9hDHKmIO86pmyfvDKAon/yNZY5b
ioptx6uSZ0RHFlCsO9eYTNeGf0CQLd1hQ+ZvaKQlEIU/BOzqcZmGWPqVGcrkZkWe
7YAnMC7VmWQxDH/jLsfhyNg2fZuvAUgKOx1jDgJKmMnYJzAvTZqTCabqmxQu/sm/
CMfzTXvXXLdXh3ACD+zc9iUO0X1N5XCihJkpHXSABb9Z2vYwEEAMk7c0nbYT+oZp
lTKTCl8/6XCQ540oLjcrWSqolXXgR6koRGK+/fpHusYB/IlX99mP644svWlFpLyZ
FL3FuGOVi6kXOYz9tlINsiTAYKnyu5xHksoBYOcUxes5SziMJOtoolre3I8aqq+7
JAVFU5Bq0nwrXBSv9vxRDNDXeNNpUCDF5YRn3CJgCxyFV/S0jGKxUpqBSiVfnOJp
aFpPXWDV5wD1ZulGSO5nRXa/AmvBabL9XDlqs2xL27WjuJtq5H1HAr2NLn1/NilJ
nF0obZuR+x7H50wXUcW2mwGl7YEUQwKnkhU6HwXCkP5QYaw5bxrBYmL/kSSVb8vc
OX7rmsJBENBfs0ooq4J09R7deSlxcMFwVM25aiVo7IaYGNqgWhKL1dWXwqhlzR2E
ft8Xi1xXFO6z4j3Zw1oWQptLMx7wjZZlLby/wW2xz2uS7K3UzQ9UMaSHRCzu4wR2
TSh5RVw1HvlBo1xCr1fIcAHypdxfxvhkD3KIsyo69X9LAlfFIv4w2afotXrQaeHi
81yzgMgpNUYKHC8/BwVJjDXHO+5E5MbRx5yfDp4E4sZGFXiQVRCH4OI5bC+oCOPx
mcg4rli5CAtuIkZ2RWbGZGpX82NXtb8nKTPqdSpEoJaljogkJYcqvY0D5rLlFewt
TfTALPIGlY7LN9h3x7YDHfPtMF97TXXDlbBNMcJVuWl8GYo7C77GJ/fkpjqOcDuN
+5Uv3o0ozDySyiCzPqa7YcAEDmKxFVvQ8jr7lD7zWRhXSNdgXniYC7GO2YAcILJa
ZmzO9terrejN4t3tJgicyVSOHtrBotfJeJnSMZwV+AL5U1gmltYaXLKuPoYerxWl
18kWksiclmiuIwCb22ChB8LSTJTrHih5sUI9i//BCYWHKRUhMKuD/JBhAc4zWvp4
5cxjYvkp4VMeAMDZ1mzaylFk9AqN9rvMad9DZXF5RcrrcW11RopwJrIL9baTUYIh
fukg6oTeRN/0QXiytcCvblz/Pao1zyX4ffNRLN147ECZ3To346D4mOwDUI99ausP
aQT8oMrhMW3bcOE0TxQOYSZz2bwIYiE4rUjbIbai/bo5KXJzVMD5U4ZlkDj7t4Hl
PJerNpqrFzgfVEibnCBtmOfEMBAQlAE1HSH+S8CUhAhDrNzsXkDIH+kyIzBw9r0b
Va4F/XIqHVcUxbDMK4eX92JK/O8nU9/upaLR3jQEgFDUcc0JZpV5OGnQwu4xB6Vm
A0dv0M8IIJAzSym8HeOM7li1mdIi4LttfRTIehk4jYckXVdB42MEwbf27YOcmshN
Hn9AIz0oUTiprvaVeY8CYmQaquLmmBrapHYvgZkVLDXyZoiDuojBjzppgkefzr3p
rqJHqMg6HFohhUEzFXYW1VUVqnxGUj4EAaZRe59bh1q5Ed0ndM4raCJCi44TgXs3
9n3mi6kT05EXJMzrB/I9fd6iy5HMee4hE8CLugZnsgSbB9pXM4rY0I28sBNfIL2M
KDX8aOccF1MNEI/z7EZplsT2aVJMeTdoKWqvyONhD+O4LT+HyyCFDjBxcY+r/pQC
s0K6anw/EYPnzeJgB90DiDiB5+CynRAvFPVtGj4niuPxTSfsObCYM2ZYtWALWoDQ
ch6qYL8tKuxhsM9LPLaTYwlXQ3FDKpgxRNl87WE67IAVeW3YV2MW+Q0HdHfIDkTb
29Bey5BdcPB+w5HiRPxUYysZMnLKDMhqzzJTJxO+CXIAV30CZdtZ9pLkZRpIMJ+f
ZK5nlvmzONmgrgrhV7BISenyIZ/gdpu/Pdp+11bZkddB0ly0aP0XlrDYmAiKhJNI
rgFKIbuxh2e8js/4uzkhCVuCySsdB+GBG2bfnJjvNdNmTS0XF/BFjt//oJptqVD+
B6tVoSsavn3QHeYDNqSkGhqt2Jx8WxpVowPOXdx4pg25jHnCuqgO4yZs0lCso55w
jCDLU7gt/+PAP6k//cjMO8DKBCh7EKSx0cMYusQEnk3z/FLUMalWrx69jG26pdxQ
khaRK67z9LoDnqOOf7cHKSDKSk7Zql9Ze2WQbB9Ev+Jr4Bjp+5fts2vizDiiTq34
VouUzl+B76yPo47pychQ1I7QBkB9hQ+oDF4Tk5AXBLD+LI8DUMMrX2smpzSPPm1X
NoQWcu63ARsXX3PbhilQZg6ck+M6ofDH8dE/oUTusZJwS3y8dT9VGonCty+Tbfx4
4U8vVMBN5wveE3P7KlwaDDcEQuoWk2agzNBNkA8E4Lolsgm6SJNv4as+skDJSlpT
IIl1lFkwjUruTYLb7XBd8cHqfFmgjAf4Wzcd1M9oGkUGhm+mz2aS6/K0p5GRdtWb
6oV88zdU2y3QYlSkgh+9xiDsTSIl4dgTTm7ieXedQ4M/RSk1bB1oguE6go5REe4J
DO3ORmozAoRDKEE299NaT1XoAQbEjzBfhnqc71VkLvX2jRdAZgpcmT4zUhFY+ene
uRpwKicrXkqLzm+KHixhf5BMHvmJbhQmEjlI5cNtLG1cPdkUUfU5Dw9uzBAmtD7/
rhi4xLW4xEQz08x2HvyuCgaByvr+1soD1E0v7t3MSyVRY7dFUIQkrpH6xlXwtHCm
+3nox0Kd/8RRmcwt+yRUPjBJlvzKvGYWqS+JvSfXDb+v9D4g6rawln7MlVRgVVFM
WpZZAiVq3HQjM5A/fszJQI8GaB92X5LlSAg/IvAT9J/DOdGxwZ8FFlKLY20ZtbHC
aLhVsueU3r/cL9FoR3FA4eP2oDL36JJwEqy05Hpm6ZQI1Mw3Ylf6BPm2W2ZoYH/K
9oHGRpojzdnLVDQxszMF0oHv6ymWDRfUmq5IhCvNI6YiFb0bv/r6tMq2irBpxQ7a
V1LUS3AXkDhPcGntPN7SPIaP0uKUUh6fl+VPkFVlJbiSBv23R2AzSW/RgC3LHWqS
DJjga7tj4FHa5C71R8OwiddR0D4sCbe6YQcmecQbEtez+lsp/P44/2yTrh2Dzruh
2AypzQXdZjVWsyqNRGK/eCURhNy7RqF4qnPXZiH1ZXVSYF9HP0pePP8mumK2bHrM
V7hOzX9+hKOuvwv4QAJgYoN8gUmQ+fRRElM17SJG+JPlNYDrmmw4rKwfxdN2DUnN
rI0J84Qh7TMLSIFtyhWgur6IKvcYLWTVW6vOsGWNV7iBAfD+WsXDERTLu7aCiQh0
a2bZ0HeonuBkEtSi1RwsDhrd9D97fMJu4jH11v3bawBv2CewuC5ev/hi8yJCZR+G
AWe+ELIhMOdbQSOQOSpvxXSXOc8LOA4hZPHy7xG0Ioj+YkSqitdJ/CVBh5yKJNzR
TDzmQOALTd5DbLF4YBl0jUs3kxT4VNijg2IhdKBme93Q9LE+hkrLN7YOnFW3shDO
cY7s5SGxRYHjWFERSd9T/cReuJFNwzUbDxtTVUqT9g9LT/kUzTMfaVY/TmPvcxnu
5VBaUdycTMb0ooj16/XuBqn8M+uaMTZzLSwZBVlDrMHrq1SCaLtxuppksbWI5+im
tyI0eKpsv3YQNi7439NEY5Vx2IZuBW+MoaMbh6m7OWplbJzO9ek4TeV0GqVmzJmZ
b5GeAUJ4mgUpqWGRszziRHb+4fk0QtAbk06amZXgQDWw8nl9LbziWBvWAZTUID01
WwXGYrueGy4ILPQsAUQBI0YTF4P+FHeDqmL9wfcmejfotAJToIxURoUNLQc9p9cG
Z/kP547emNN9nHUkuJMWSNqphraeEHXZOYVOl76hirYzIfxES6jBV9hJw4HallAJ
vjENgrWmA4UjIesO43BXi5skc//RNnQ8ZsvWYTY5EJDCAh41JNIQD2RR694jA9wT
7IwSlQA5J6LekUf+q6nG0rnJH0A56qOasyeD2Tu4vvrPz9l2lY7aZ5NxHQPx0UP7
oontpUdJcBpcYpMpYcK0enstOqwCHudWUlNvEVsLzquAIZW1oGQ9eKAi4E0HZday
EeuNyu47EKmKQAeCnN2gzMixYERyyBTSvkWVBN8x0V3da1qulPzM+WqekkoEUtlt
LHPRl4QM0HZgZRQ8YnUecV0QOeLl13EjZpgXtkyf1pcxN/aL+nd6YVEnZvSKglfG
nfJ36OJE2oDaksTY1ddr/r3I/9EYLbwGKOjOn9rWlGvjryQJeWpnY79lt4Js52PN
CzmWtEYtVdSCmcSOzbKPqOZxn08O65uel8THk+ZDElGMAvtj9MDPHRHchpZb1dS7
+9p5iwaRQb3BcWqVcoAu3bW7T3K/PDva5+45Kh7FSJXJZyBeI0gKHTnAXDQo0dkG
BhFcrN/t+kJbkav1U7clrg1Kv9vwOYcqfz7oUxUTrUQpcSi1AlQ4X7UZrMk3KlD5
GQhiCb+3SxY7DriyCvMkki+sWB0km4doNjpAPIP1t0MH9YSqYLouSH8vyWK7bHW8
jkUyEdXWnyd52lO1yNYuydTODfNr8YEKC0jYk/TZLdBuQ1F0Uz/CY+dlriCd0p09
7hEEXVxy/b6eQYZv5U8XTB4UWaQHWs5cE4eh6t+PV3lq6K3e3aHjsQDtPD6k7u7z
tIHMATE8ZLujJSd9m8FVo7cIvF1RLtDssM2hW9wyBRuX5UCQ0WH4VGy5mHwwU5V6
Cc9T2EHqACKyrExaxqHvHUaJn6Iv16WUif61Cew1ZjSpaOLoVD/YRJBmVkylJzvS
zMLbfYtwB/sTnJ0wtM2xlhGGE8dtJl87ES4jprahajJk3dmbpudIpBVrTs3XrNI0
LLP7+Pp0JOpmeVbtsgD6Eqp9t2BdRgdr67JC0KChfBvC197hkEdp2NJ2Fo6ixYVI
+o29Uj5Iw79mN8NHDImaOyYsr7/cSv2eQ0bRP0kYphXYi2BCE1gdUwiewYEXDa5+
D2qNXZDeAdLe2SckiyHdhluCeheHg4Ctec/CCmAEV52exdmMfHbDDsL5mr0UdpuB
`protect end_protected
