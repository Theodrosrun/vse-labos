/*******************************************************************************
HEIG-VD
Haute Ecole d'Ingenerie et de Gestion du Canton de Vaud
School of Engineering and Management Vaud
********************************************************************************
REDS Institute
Reconfigurable and Embedded Digital Systems
********************************************************************************

File     : min_max_top_tb.sv
Author   : Yann Thoma
Date     : 07.10.2024

Context  : min max component testbench

********************************************************************************
Description : This testbench is decomposed into stimuli
              generation and verification, with the use of interfaces.

********************************************************************************
Dependencies : -

********************************************************************************
Modifications :
Ver   Date        Person     Comments
1.0   07.10.2024  TMU        Initial version

*******************************************************************************/

interface min_max_in_itf#(int VALSIZE);
    logic[1:0] com;
    logic[VALSIZE-1:0] max;
    logic[VALSIZE-1:0] min;
    logic osci;
    logic[VALSIZE-1:0] value;
endinterface

interface min_max_out_itf#(int VALSIZE);
    logic[2**VALSIZE-1:0] leds;
endinterface

module min_max_top_tb#(int VALSIZE, int TESTCASE, int ERRNO);

    timeunit 1ns;         // Definition of the time unit
    timeprecision 1ns;    // Definition of the time precision
   
    // Reference
    logic[2**VALSIZE-1:0] leds_ref;
   
    // Timings definitions
    time sim_step = 10ns;
    time pulse = 0ns;
    logic synchro = 0;
   
    always #(sim_step/2) synchro = ~synchro;
   
    // Interfaces
    min_max_in_itf input_itf();
    min_max_out_itf output_itf();

    // Erros values
    logic error_signal = 0;
    int nb_errors = 0;

    // Typedef
    typedef logic[VALSIZE-1:0] input_t;
    typedef logic[2**VALSIZE-1:0] output_t;

    // DUV instantiation
    min_max_top#(VALSIZE, ERRNO) duv(.com_i(input_itf.com),
                                     .max_i(input_itf.max),
                                     .min_i(input_itf.min),
                                     .osc_i(input_itf.osci),
                                     .val_i(input_itf.value),
                                     .leds_o(output_itf.leds));

    // ***********************************************
    // ******************** class ********************
    // ***********************************************

    class RBase;
        rand logic[1:0] com;
        rand input_t max;
        rand input_t min;
        rand logic osci;
        rand input_t value;

        constraint max_bigger_than_min {
            max > min;
        }
    endclass

    class RCoverage extends RBase;
        covergroup cg;
            option.at_least = 1000;

            coverpoint com { 
                bins values[] = {0, 1, 2, 3};
            }

            coverpoint max { 
                bins values[VALSIZE] = {[0:2**VALSIZE-1]};
            }

            coverpoint min { 
                bins values[VALSIZE] = {[0:2**VALSIZE-1]};
            }

            coverpoint osci { 
                bins values = {0,1};
            }

            coverpoint value { 
                bins values[VALSIZE] = {[0:2**VALSIZE-1]};
            }
        endgroup

        function new();
            cg = new();
        endfunction

        task start();
            automatic int generation_count = 0;
            while (cg.get_coverage() < 100) begin
                generation_count++;
                if (!randomize()) begin
                    $display("%m: randomization failed");
                end else begin
                    input_itf.com = this.com;
                    input_itf.max = this.max;
                    input_itf.min = this.min;
                    input_itf.osci = this.osci;
                    input_itf.value = this.value;
                    @(posedge(synchro));
                    cg.sample();
                    $display("coverage rate: %0.2f%%", cg.get_coverage());
                end
            end
            $display("coveraged finished\n");
        endtask
    endclass

    class RTest extends RBase;
        task start();
            automatic int generation_count = 0;

            for(integer i = 0; i < 1000; i++)begin
                generation_count++;
                if (!randomize()) begin
                    $display("%m: randomization failed");
                end else begin
                    input_itf.com = this.com;
                    input_itf.max = this.max;
                    input_itf.min = this.min;
                    input_itf.osci = this.osci;
                    input_itf.value = this.value;
                    @(posedge(synchro));
                end
            end
            $display("randomization finished\n");
        endtask
    endclass

    class RTestOutOfRangeMin extends RTest;
        constraint value_smaller_than_min {
            value < min;
        }
    endclass

    class RTestOutOfRangeMax extends RTest;
        constraint value_bigger_than_max {
            value > max;
        }
    endclass
    
    class RTestBoundariesMin extends RTest;
        constraint boundaries {
            value == min;
        }
    endclass

    class RTestBoundariesMax extends RTest;
        constraint boundaries {
            value == max;
        }
    endclass

    task test_coverage();
        automatic RCoverage rt = new();
        rt.start();
    endtask

    task test_randomized_out_of_range_min();
        automatic RTestOutOfRangeMin rt = new();
        rt.start();
    endtask

    task test_randomized_out_of_range_max();
        automatic RTestOutOfRangeMax rt = new();
        rt.start();
    endtask

    task test_randomized_boundaries_min();
        automatic RTestBoundariesMin rt = new();
        rt.start();
    endtask

    task test_randomized_boundaries_max();
        automatic RTestBoundariesMax rt = new();
        rt.start();
    endtask

    task test_value_equals_max();
        input_itf.min = 0;
        input_itf.max = 2**VALSIZE - 1;
        input_itf.value = 2**VALSIZE - 1;
        input_itf.com = 2'b00;
        input_itf.osci = 0;
        @(posedge(synchro));
    endtask

    task test_osci();
        input_itf.min = 5;
        input_itf.max = 10;
        input_itf.value = 7;
        input_itf.com = 2'b00;
        input_itf.osci = 1'b0;
        @(posedge(synchro));

        assert (output_itf.leds[10:8] == 3'b000) else $display("%m: LEDs should be off");
        input_itf.osci = 1'b1;  
        @(posedge(synchro));

        assert (output_itf.leds[10:8] == 3'b111) else $display("%m: LEDs should be on with low intensity");
        input_itf.osci = 1'b0;
        @(posedge(synchro));

        assert (output_itf.leds[10:8] == 3'b000) else $display("%m: LEDs should be off again");
    endtask

    // ***********************************************
    // ******************* Program *******************
    // ***********************************************

    task tests(int TESTCASE);
        if (TESTCASE == 0) begin
            $display("Running all test scenarios...");
            test_coverage();
            test_randomized_out_of_range_min();
            test_randomized_out_of_range_max();
            test_randomized_boundaries_min();
            test_randomized_boundaries_max();
            test_value_equals_max();
            test_osci();
        end
        else begin
            case(TESTCASE)
                1: test_coverage();
                2: test_randomized_out_of_range_min();
                3: test_randomized_out_of_range_max();
                4: test_randomized_boundaries_min();
                5: test_randomized_boundaries_max();
                6: test_value_equals_max();
                7: test_osci();
                default: begin
                    $display("Invalid TESTCASE: %d", TESTCASE);
                    $finish;
                end
            endcase
        end
    endtask

    task compute_reference(logic[1:0] com, input_t min, input_t max, input_t value, logic osci, output output_t leds);
        leds = {2**VALSIZE{1'b0}};
        
        case (com)
            2'b00: // Normal mode
            begin 
                if (value >= min && value <= max) begin
                    for (integer i = min; i <= value; i++) begin
                        leds[i] = 1;
                    end
                    for (integer i = value + 1; i <= max; i++) begin
                        leds[i] = osci;
                    end
                end
            end
            
            2'b01: // Linear mode
            begin
                for (integer i = 0; i <= value; i++) begin
                    leds[i] = 1;
                end
            end

            2'b10: // Test all OFF 
            begin
                // Set to 0 by default
            end

            2'b11: // Test all ON
            begin
                leds = {2**VALSIZE{1'b1}}; 
            end
        endcase
    endtask

    task compute_reference_task;
        forever begin
            @(posedge(synchro));
            #1;
            compute_reference(input_itf.com, input_itf.min, input_itf.max, input_itf.value, input_itf.osci, leds_ref);
        end
    endtask

    task verification;
        @(negedge(synchro));
        forever begin
            if (output_itf.leds !== leds_ref) begin
                nb_errors++;
                $error("%m: Error for com = %b, min = %d, max = %d, value = %d \nExpected: %b \nObserved: %b", 
                       input_itf.com, input_itf.min, input_itf.max, input_itf.value, leds_ref, output_itf.leds);
                error_signal = 1;
                #pulse;
                error_signal = 0;
            end
            @(negedge(synchro));
        end
    endtask

    initial begin
        $display("\nStarting simulation");
        fork
            tests(TESTCASE);
            compute_reference_task;
            verification;
        join_any

        if (nb_errors > 0)
            $display("Number of errors : %d", nb_errors);
        else
            $display("No errors");

        $display("Simulation finished\n");
        $finish;
    end

endmodule
