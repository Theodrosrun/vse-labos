`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
TwAUF6h1pxEsJN/pD6+S7GkfxnvFy1vtiYUwQQp8WT21Mpmbn/7TU//YCEboIHqC
JSsxJ3cYTNJbZeY1vIm/b1dJHNu2WuJwObJwbAkxz5HcNLnBXDY957g/u0DSaGFu
CO+Rw2xv2xR4g9NPPaTFZLeP7Q6JAuTHC4mZP9LXouZ6QDRtTW21DGl4gmB0sXtV
iKnhMnO28YpkVJQGvm/7wmdqX5hRbTA8d3BTjmnhZCozgekZ0saDY5rqrRl4NMOo
RRtJSbEZi4mTJJINHeQmXnUijaSFOH0QyApiqZf48jjutngq4c2cMbhruEagr77R
5wkwx1/D9U6iKCHerWUOxA==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1520 )
`protect data_block
ZK9djo00ag4nXK6qc1p5Mw3hF+9R7wa7ch/mjsGTOlhFpK8iIz6K1RWk6VifZoz+
6P4FssrG7QEndroglXVYuSqyh5ZlqdwqQQPWpZjeEsU2r57+Y5ruk/CUhMnYVW4C
Ncw6pp6krV0Hp7rkuEiuGfs69hAcW0klwniVV/FqFKvactl9Zy0fJ5qR3cuOTmmf
ZT7Vb7zdtT337wGepizc20gxABY8cPO6iLyfS04uOapdAmIX2cN3S6Y0NVsBKVR4
Z8c0PuvEURn0Z3uohWMqKC+QvZaaDZuPtKZVvbjrlI7p45kp8CMHtm7+TljqpVIm
KilCrPHxynM36fPRKAusAliqk0PLyHRty+LICKVo08V9p78AlFkEtK/WiVY9ZKO2
0jMuWWsve8J+utAa9VRi1jEaK1bl/4q0jf7fO7MRROu4bNlH9j6A2IaUvznkypM1
zTKOxwG5dG6zlnhlJj3fvBQVop7XwwB9TZcJ5x4kxrHnj3sRDen1MY1QZX/wuFLs
VOqK5D2qbR3d41kqg5mkmiarN3mwtP4nb04Z4/maOwkfPKFCwPGeXJTOUz5JIV2i
cQZSKUI4asXCbqwOjwqXwgqgAavmLVMP8aZKfYpmUiAsT68n/8x+1AdHSPOqXWTG
CiSGxiWuB7SMgx9ZTknn3B35MEfsPRIPd7GNOwJQaTbVrWBklHLdnrllKpFw3BAG
HbD5PSZHtqpJbhjTY68tnx0EydoAMf0jazYrUcKgwrQONwYLRD/ZLr/n1QNnela1
UekDZb80Fny9sv16WGhpyTgG8QmOoCaiuOKkKS4i9hhFiT9KzbomRWWVDr87NwE5
r/gd0j80h9OPXGC4XnvnRZzxN57wQ9BgG8U9Lsi/ggJ9OTQ8a08VngWVcsmzYkoX
0MXcG6wm3GLDTa5rWo3maPoKrpGMR5ZNzKJj1ki18IxjJmLi6WCoLo8AHoQcAHHI
gvs9JiKDCHebWbXZQeVrAAh+5TV0FuayrmZ/b8jP1/fMQ5mSp+hzv0cvO1iUdv3s
+kUjgpqQlKzNsgGYRJPYIwE7QuQM5UB38+LTX3yGtjQpGcTJo2lWtgsgrPbpMDsA
8ATLm/LFZ3OdXX4YEXjEkTqXQYc+WGnj7ReZNldjjbblzJRab/3g/x6a0mJ/vZAH
6pXHw8LJdLQ+gR+O8O62lyUTc2LNr0lOVJd8XQS6l4WV+Hp7lRwW5CH1d0rESIue
NOl1Xc5sOLc0akxbbCYcP+8Ay+WllVlBReLBY6X2rpZS1QFJTEFMPdxY0D95Hs/0
+KuVUswD0i3FQTyv28Jm+jFTpHS+WRWH9tM5l1D/KJgm2Nqvkr9ZqNR5ZclgpOS+
uHamorF7Gpo96suGvnCBJfatBVpqaS5If1ZjYHewfvx6r/TSRMmCXVRUYCDjXSJg
XcnMvRmIZrIMaig9/TZs9lB9O8HLKO4c3qJLG1mRjfsWl6kD2xWBmsnY+yqjyWIO
7SROOTrUvKjSYKHFnNreLYflD1ctPYq0NvY64hteIMW6gSq1uTvGfvJ6P68LFWWA
9iYXGDc6FUuAmIIYVb4AjJ0aRYP5mAnd/2BIXzQ8hQ0t8P4p4TA4WhWiOsTH7NNa
8ecMTNjoR5gfGH/p2Ny7fwcH12H3yCHcvkCzt8OJq/ycAM7/9JGf9qfoympHe+7Y
Wgb5OYbwPZLoF/5elzJIkbBYuBnPJlMn5H2Tgk5U1yDpJ5PluDQwd2DYJRBVmMa4
Joohm5HbZ126orkAGcD0ez51+w9W9sOc2UnhYOpgUBM/UR2GOa4LNsDMSzDu/Yqt
lxwGoenUxK4X7IgZUYaORsTRJSJ6fSsJHUZN+uyKPq2TEE2HI7rIkxnasUFgZ3ip
HWvJ+H8UoNqPmXv0vJMDwppudF2Asewnh6T5MR5s7w7IcRe6Oj84F/0yD7KSH3pP
6ZAYrUVQJOucP470HuxxK2SrrPBxdIjEdPCZm9wJJ86Pf3hd1FsjPFEJQpBHVui7
Xu5pjpbYEslFZaDkUc2A76pC4r/wjOzCAjwCIuqqWkk=
`protect end_protected
